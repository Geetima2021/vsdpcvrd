module rvmyth (clk,
    reset,
    VPWR,
    VGND,
    out);
 input clk;
 input reset;
 input VPWR;
 input VGND;
 output [7:0] out;

 sky130_fd_sc_hd__inv_2 _09635_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .Y(_04646_));
 sky130_fd_sc_hd__buf_2 _09636_ (.A(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__nand2_4 _09637_ (.A(CPU_is_s_instr_a4),
    .B(CPU_valid_a4),
    .Y(_04648_));
 sky130_fd_sc_hd__buf_2 _09638_ (.A(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__buf_2 _09639_ (.A(\CPU_dmem_addr_a4[1] ),
    .X(_04650_));
 sky130_fd_sc_hd__buf_2 _09640_ (.A(\CPU_dmem_addr_a4[0] ),
    .X(_04651_));
 sky130_fd_sc_hd__buf_2 _09641_ (.A(\CPU_dmem_addr_a4[3] ),
    .X(_04652_));
 sky130_fd_sc_hd__buf_2 _09642_ (.A(\CPU_dmem_addr_a4[2] ),
    .X(_04653_));
 sky130_fd_sc_hd__or4_4 _09643_ (.A(_04650_),
    .B(_04651_),
    .C(_04652_),
    .D(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__buf_2 _09644_ (.A(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__nor2_4 _09645_ (.A(_04649_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__buf_2 _09646_ (.A(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__buf_2 _09647_ (.A(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__buf_2 _09648_ (.A(CPU_reset_a4),
    .X(_04659_));
 sky130_fd_sc_hd__buf_2 _09649_ (.A(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__buf_2 _09650_ (.A(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__buf_2 _09651_ (.A(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__buf_2 _09652_ (.A(_04656_),
    .X(_04663_));
 sky130_fd_sc_hd__buf_2 _09653_ (.A(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__nor2_4 _09654_ (.A(\CPU_Dmem_value_a5[0][30] ),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a211o_4 _09655_ (.A1(_04647_),
    .A2(_04658_),
    .B1(_04662_),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__inv_2 _09656_ (.A(_04666_),
    .Y(_01548_));
 sky130_fd_sc_hd__inv_2 _09657_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .Y(_04667_));
 sky130_fd_sc_hd__buf_2 _09658_ (.A(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__nor2_4 _09659_ (.A(\CPU_Dmem_value_a5[0][29] ),
    .B(_04664_),
    .Y(_04669_));
 sky130_fd_sc_hd__a211o_4 _09660_ (.A1(_04668_),
    .A2(_04658_),
    .B1(_04662_),
    .C1(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__inv_2 _09661_ (.A(_04670_),
    .Y(_01547_));
 sky130_fd_sc_hd__inv_2 _09662_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .Y(_04671_));
 sky130_fd_sc_hd__buf_2 _09663_ (.A(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__nor2_4 _09664_ (.A(\CPU_Dmem_value_a5[0][28] ),
    .B(_04664_),
    .Y(_04673_));
 sky130_fd_sc_hd__a211o_4 _09665_ (.A1(_04672_),
    .A2(_04658_),
    .B1(_04662_),
    .C1(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__inv_2 _09666_ (.A(_04674_),
    .Y(_01546_));
 sky130_fd_sc_hd__inv_2 _09667_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .Y(_04675_));
 sky130_fd_sc_hd__buf_2 _09668_ (.A(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_4 _09669_ (.A(\CPU_Dmem_value_a5[0][27] ),
    .B(_04664_),
    .Y(_04677_));
 sky130_fd_sc_hd__a211o_4 _09670_ (.A1(_04676_),
    .A2(_04658_),
    .B1(_04662_),
    .C1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__inv_2 _09671_ (.A(_04678_),
    .Y(_01545_));
 sky130_fd_sc_hd__inv_2 _09672_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .Y(_04679_));
 sky130_fd_sc_hd__buf_2 _09673_ (.A(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__buf_2 _09674_ (.A(_04661_),
    .X(_04681_));
 sky130_fd_sc_hd__buf_2 _09675_ (.A(_04663_),
    .X(_04682_));
 sky130_fd_sc_hd__nor2_4 _09676_ (.A(\CPU_Dmem_value_a5[0][26] ),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__a211o_4 _09677_ (.A1(_04680_),
    .A2(_04658_),
    .B1(_04681_),
    .C1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__inv_2 _09678_ (.A(_04684_),
    .Y(_01544_));
 sky130_fd_sc_hd__inv_2 _09679_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .Y(_04685_));
 sky130_fd_sc_hd__buf_2 _09680_ (.A(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__nor2_4 _09681_ (.A(\CPU_Dmem_value_a5[0][25] ),
    .B(_04682_),
    .Y(_04687_));
 sky130_fd_sc_hd__a211o_4 _09682_ (.A1(_04686_),
    .A2(_04658_),
    .B1(_04681_),
    .C1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__inv_2 _09683_ (.A(_04688_),
    .Y(_01543_));
 sky130_fd_sc_hd__inv_2 _09684_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .Y(_04689_));
 sky130_fd_sc_hd__buf_2 _09685_ (.A(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__buf_2 _09686_ (.A(_04657_),
    .X(_04691_));
 sky130_fd_sc_hd__nor2_4 _09687_ (.A(\CPU_Dmem_value_a5[0][24] ),
    .B(_04682_),
    .Y(_04692_));
 sky130_fd_sc_hd__a211o_4 _09688_ (.A1(_04690_),
    .A2(_04691_),
    .B1(_04681_),
    .C1(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__inv_2 _09689_ (.A(_04693_),
    .Y(_01542_));
 sky130_fd_sc_hd__inv_2 _09690_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .Y(_04694_));
 sky130_fd_sc_hd__buf_2 _09691_ (.A(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__nor2_4 _09692_ (.A(\CPU_Dmem_value_a5[0][23] ),
    .B(_04682_),
    .Y(_04696_));
 sky130_fd_sc_hd__a211o_4 _09693_ (.A1(_04695_),
    .A2(_04691_),
    .B1(_04681_),
    .C1(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__inv_2 _09694_ (.A(_04697_),
    .Y(_01541_));
 sky130_fd_sc_hd__inv_2 _09695_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .Y(_04698_));
 sky130_fd_sc_hd__buf_2 _09696_ (.A(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__nor2_4 _09697_ (.A(\CPU_Dmem_value_a5[0][22] ),
    .B(_04682_),
    .Y(_04700_));
 sky130_fd_sc_hd__a211o_4 _09698_ (.A1(_04699_),
    .A2(_04691_),
    .B1(_04681_),
    .C1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__inv_2 _09699_ (.A(_04701_),
    .Y(_01540_));
 sky130_fd_sc_hd__inv_2 _09700_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .Y(_04702_));
 sky130_fd_sc_hd__buf_2 _09701_ (.A(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__nor2_4 _09702_ (.A(\CPU_Dmem_value_a5[0][21] ),
    .B(_04682_),
    .Y(_04704_));
 sky130_fd_sc_hd__a211o_4 _09703_ (.A1(_04703_),
    .A2(_04691_),
    .B1(_04681_),
    .C1(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__inv_2 _09704_ (.A(_04705_),
    .Y(_01539_));
 sky130_fd_sc_hd__inv_2 _09705_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .Y(_04706_));
 sky130_fd_sc_hd__buf_2 _09706_ (.A(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__buf_2 _09707_ (.A(_04661_),
    .X(_04708_));
 sky130_fd_sc_hd__buf_2 _09708_ (.A(_04663_),
    .X(_04709_));
 sky130_fd_sc_hd__nor2_4 _09709_ (.A(\CPU_Dmem_value_a5[0][20] ),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__a211o_4 _09710_ (.A1(_04707_),
    .A2(_04691_),
    .B1(_04708_),
    .C1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__inv_2 _09711_ (.A(_04711_),
    .Y(_01538_));
 sky130_fd_sc_hd__inv_2 _09712_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .Y(_04712_));
 sky130_fd_sc_hd__buf_2 _09713_ (.A(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__nor2_4 _09714_ (.A(\CPU_Dmem_value_a5[0][19] ),
    .B(_04709_),
    .Y(_04714_));
 sky130_fd_sc_hd__a211o_4 _09715_ (.A1(_04713_),
    .A2(_04691_),
    .B1(_04708_),
    .C1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__inv_2 _09716_ (.A(_04715_),
    .Y(_01537_));
 sky130_fd_sc_hd__inv_2 _09717_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .Y(_04716_));
 sky130_fd_sc_hd__buf_2 _09718_ (.A(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__buf_2 _09719_ (.A(_04663_),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_4 _09720_ (.A(\CPU_Dmem_value_a5[0][18] ),
    .B(_04709_),
    .Y(_04719_));
 sky130_fd_sc_hd__a211o_4 _09721_ (.A1(_04717_),
    .A2(_04718_),
    .B1(_04708_),
    .C1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__inv_2 _09722_ (.A(_04720_),
    .Y(_01536_));
 sky130_fd_sc_hd__inv_2 _09723_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .Y(_04721_));
 sky130_fd_sc_hd__buf_2 _09724_ (.A(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__nor2_4 _09725_ (.A(\CPU_Dmem_value_a5[0][17] ),
    .B(_04709_),
    .Y(_04723_));
 sky130_fd_sc_hd__a211o_4 _09726_ (.A1(_04722_),
    .A2(_04718_),
    .B1(_04708_),
    .C1(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__inv_2 _09727_ (.A(_04724_),
    .Y(_01535_));
 sky130_fd_sc_hd__inv_2 _09728_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .Y(_04725_));
 sky130_fd_sc_hd__buf_2 _09729_ (.A(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__nor2_4 _09730_ (.A(\CPU_Dmem_value_a5[0][16] ),
    .B(_04709_),
    .Y(_04727_));
 sky130_fd_sc_hd__a211o_4 _09731_ (.A1(_04726_),
    .A2(_04718_),
    .B1(_04708_),
    .C1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__inv_2 _09732_ (.A(_04728_),
    .Y(_01534_));
 sky130_fd_sc_hd__inv_2 _09733_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .Y(_04729_));
 sky130_fd_sc_hd__buf_2 _09734_ (.A(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_4 _09735_ (.A(\CPU_Dmem_value_a5[0][15] ),
    .B(_04709_),
    .Y(_04731_));
 sky130_fd_sc_hd__a211o_4 _09736_ (.A1(_04730_),
    .A2(_04718_),
    .B1(_04708_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__inv_2 _09737_ (.A(_04732_),
    .Y(_01533_));
 sky130_fd_sc_hd__inv_2 _09738_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .Y(_04733_));
 sky130_fd_sc_hd__buf_2 _09739_ (.A(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__buf_2 _09740_ (.A(_04661_),
    .X(_04735_));
 sky130_fd_sc_hd__buf_2 _09741_ (.A(_04656_),
    .X(_04736_));
 sky130_fd_sc_hd__nor2_4 _09742_ (.A(\CPU_Dmem_value_a5[0][14] ),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__a211o_4 _09743_ (.A1(_04734_),
    .A2(_04718_),
    .B1(_04735_),
    .C1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__inv_2 _09744_ (.A(_04738_),
    .Y(_01532_));
 sky130_fd_sc_hd__inv_2 _09745_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .Y(_04739_));
 sky130_fd_sc_hd__buf_2 _09746_ (.A(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__nor2_4 _09747_ (.A(\CPU_Dmem_value_a5[0][13] ),
    .B(_04736_),
    .Y(_04741_));
 sky130_fd_sc_hd__a211o_4 _09748_ (.A1(_04740_),
    .A2(_04718_),
    .B1(_04735_),
    .C1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__inv_2 _09749_ (.A(_04742_),
    .Y(_01531_));
 sky130_fd_sc_hd__inv_2 _09750_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .Y(_04743_));
 sky130_fd_sc_hd__buf_2 _09751_ (.A(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__buf_2 _09752_ (.A(_04663_),
    .X(_04745_));
 sky130_fd_sc_hd__nor2_4 _09753_ (.A(\CPU_Dmem_value_a5[0][12] ),
    .B(_04736_),
    .Y(_04746_));
 sky130_fd_sc_hd__a211o_4 _09754_ (.A1(_04744_),
    .A2(_04745_),
    .B1(_04735_),
    .C1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__inv_2 _09755_ (.A(_04747_),
    .Y(_01530_));
 sky130_fd_sc_hd__inv_2 _09756_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .Y(_04748_));
 sky130_fd_sc_hd__buf_2 _09757_ (.A(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_4 _09758_ (.A(\CPU_Dmem_value_a5[0][11] ),
    .B(_04736_),
    .Y(_04750_));
 sky130_fd_sc_hd__a211o_4 _09759_ (.A1(_04749_),
    .A2(_04745_),
    .B1(_04735_),
    .C1(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__inv_2 _09760_ (.A(_04751_),
    .Y(_01529_));
 sky130_fd_sc_hd__inv_2 _09761_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .Y(_04752_));
 sky130_fd_sc_hd__buf_2 _09762_ (.A(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__nor2_4 _09763_ (.A(\CPU_Dmem_value_a5[0][10] ),
    .B(_04736_),
    .Y(_04754_));
 sky130_fd_sc_hd__a211o_4 _09764_ (.A1(_04753_),
    .A2(_04745_),
    .B1(_04735_),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__inv_2 _09765_ (.A(_04755_),
    .Y(_01528_));
 sky130_fd_sc_hd__inv_2 _09766_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .Y(_04756_));
 sky130_fd_sc_hd__buf_2 _09767_ (.A(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__nor2_4 _09768_ (.A(\CPU_Dmem_value_a5[0][9] ),
    .B(_04736_),
    .Y(_04758_));
 sky130_fd_sc_hd__a211o_4 _09769_ (.A1(_04757_),
    .A2(_04745_),
    .B1(_04735_),
    .C1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__inv_2 _09770_ (.A(_04759_),
    .Y(_01527_));
 sky130_fd_sc_hd__inv_2 _09771_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .Y(_04760_));
 sky130_fd_sc_hd__buf_2 _09772_ (.A(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__buf_2 _09773_ (.A(_04661_),
    .X(_04762_));
 sky130_fd_sc_hd__buf_2 _09774_ (.A(_04656_),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_4 _09775_ (.A(\CPU_Dmem_value_a5[0][8] ),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__a211o_4 _09776_ (.A1(_04761_),
    .A2(_04745_),
    .B1(_04762_),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__inv_2 _09777_ (.A(_04765_),
    .Y(_01526_));
 sky130_fd_sc_hd__inv_2 _09778_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .Y(_04766_));
 sky130_fd_sc_hd__buf_2 _09779_ (.A(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__nor2_4 _09780_ (.A(\CPU_Dmem_value_a5[0][7] ),
    .B(_04763_),
    .Y(_04768_));
 sky130_fd_sc_hd__a211o_4 _09781_ (.A1(_04767_),
    .A2(_04745_),
    .B1(_04762_),
    .C1(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__inv_2 _09782_ (.A(_04769_),
    .Y(_01525_));
 sky130_fd_sc_hd__inv_2 _09783_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .Y(_04770_));
 sky130_fd_sc_hd__buf_2 _09784_ (.A(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__buf_2 _09785_ (.A(_04663_),
    .X(_04772_));
 sky130_fd_sc_hd__nor2_4 _09786_ (.A(\CPU_Dmem_value_a5[0][6] ),
    .B(_04763_),
    .Y(_04773_));
 sky130_fd_sc_hd__a211o_4 _09787_ (.A1(_04771_),
    .A2(_04772_),
    .B1(_04762_),
    .C1(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__inv_2 _09788_ (.A(_04774_),
    .Y(_01524_));
 sky130_fd_sc_hd__inv_2 _09789_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .Y(_04775_));
 sky130_fd_sc_hd__buf_2 _09790_ (.A(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_4 _09791_ (.A(\CPU_Dmem_value_a5[0][5] ),
    .B(_04763_),
    .Y(_04777_));
 sky130_fd_sc_hd__a211o_4 _09792_ (.A1(_04776_),
    .A2(_04772_),
    .B1(_04762_),
    .C1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__inv_2 _09793_ (.A(_04778_),
    .Y(_01523_));
 sky130_fd_sc_hd__inv_2 _09794_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .Y(_04779_));
 sky130_fd_sc_hd__buf_2 _09795_ (.A(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_4 _09796_ (.A(\CPU_Dmem_value_a5[0][4] ),
    .B(_04763_),
    .Y(_04781_));
 sky130_fd_sc_hd__a211o_4 _09797_ (.A1(_04780_),
    .A2(_04772_),
    .B1(_04762_),
    .C1(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__inv_2 _09798_ (.A(_04782_),
    .Y(_01522_));
 sky130_fd_sc_hd__inv_2 _09799_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .Y(_04783_));
 sky130_fd_sc_hd__buf_2 _09800_ (.A(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__nor2_4 _09801_ (.A(\CPU_Dmem_value_a5[0][3] ),
    .B(_04763_),
    .Y(_04785_));
 sky130_fd_sc_hd__a211o_4 _09802_ (.A1(_04784_),
    .A2(_04772_),
    .B1(_04762_),
    .C1(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__inv_2 _09803_ (.A(_04786_),
    .Y(_01521_));
 sky130_fd_sc_hd__inv_2 _09804_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .Y(_04787_));
 sky130_fd_sc_hd__buf_2 _09805_ (.A(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__buf_2 _09806_ (.A(_04660_),
    .X(_04789_));
 sky130_fd_sc_hd__buf_2 _09807_ (.A(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_4 _09808_ (.A(\CPU_Dmem_value_a5[0][2] ),
    .B(_04657_),
    .Y(_04791_));
 sky130_fd_sc_hd__a211o_4 _09809_ (.A1(_04788_),
    .A2(_04772_),
    .B1(_04790_),
    .C1(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__inv_2 _09810_ (.A(_04792_),
    .Y(_01520_));
 sky130_fd_sc_hd__inv_2 _09811_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .Y(_04793_));
 sky130_fd_sc_hd__buf_2 _09812_ (.A(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__nor2_4 _09813_ (.A(\CPU_Dmem_value_a5[0][1] ),
    .B(_04657_),
    .Y(_04795_));
 sky130_fd_sc_hd__a211o_4 _09814_ (.A1(_04794_),
    .A2(_04772_),
    .B1(_04790_),
    .C1(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__inv_2 _09815_ (.A(_04796_),
    .Y(_01519_));
 sky130_fd_sc_hd__inv_2 _09816_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .Y(_04797_));
 sky130_fd_sc_hd__buf_2 _09817_ (.A(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__nor2_4 _09818_ (.A(\CPU_Dmem_value_a5[0][0] ),
    .B(_04657_),
    .Y(_04799_));
 sky130_fd_sc_hd__a211o_4 _09819_ (.A1(_04798_),
    .A2(_04664_),
    .B1(_04790_),
    .C1(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__inv_2 _09820_ (.A(_04800_),
    .Y(_01518_));
 sky130_fd_sc_hd__inv_2 _09821_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .Y(_04801_));
 sky130_fd_sc_hd__buf_2 _09822_ (.A(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__inv_2 _09823_ (.A(\CPU_dmem_addr_a4[0] ),
    .Y(_04803_));
 sky130_fd_sc_hd__buf_2 _09824_ (.A(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__or4_4 _09825_ (.A(\CPU_dmem_addr_a4[3] ),
    .B(\CPU_dmem_addr_a4[2] ),
    .C(_04650_),
    .D(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__buf_2 _09826_ (.A(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__nor2_4 _09827_ (.A(_04649_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__buf_2 _09828_ (.A(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__buf_2 _09829_ (.A(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__buf_2 _09830_ (.A(_04808_),
    .X(_04810_));
 sky130_fd_sc_hd__nor2_4 _09831_ (.A(\CPU_Dmem_value_a5[1][31] ),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__a211o_4 _09832_ (.A1(_04802_),
    .A2(_04809_),
    .B1(_04790_),
    .C1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__inv_2 _09833_ (.A(_04812_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_4 _09834_ (.A(\CPU_Dmem_value_a5[1][30] ),
    .B(_04810_),
    .Y(_04813_));
 sky130_fd_sc_hd__a211o_4 _09835_ (.A1(_04647_),
    .A2(_04809_),
    .B1(_04790_),
    .C1(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__inv_2 _09836_ (.A(_04814_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_4 _09837_ (.A(\CPU_Dmem_value_a5[1][29] ),
    .B(_04810_),
    .Y(_04815_));
 sky130_fd_sc_hd__a211o_4 _09838_ (.A1(_04668_),
    .A2(_04809_),
    .B1(_04790_),
    .C1(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__inv_2 _09839_ (.A(_04816_),
    .Y(_01515_));
 sky130_fd_sc_hd__buf_2 _09840_ (.A(_04789_),
    .X(_04817_));
 sky130_fd_sc_hd__buf_2 _09841_ (.A(_04808_),
    .X(_04818_));
 sky130_fd_sc_hd__nor2_4 _09842_ (.A(\CPU_Dmem_value_a5[1][28] ),
    .B(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__a211o_4 _09843_ (.A1(_04672_),
    .A2(_04809_),
    .B1(_04817_),
    .C1(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__inv_2 _09844_ (.A(_04820_),
    .Y(_01514_));
 sky130_fd_sc_hd__buf_2 _09845_ (.A(_04807_),
    .X(_04821_));
 sky130_fd_sc_hd__buf_2 _09846_ (.A(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__nor2_4 _09847_ (.A(\CPU_Dmem_value_a5[1][27] ),
    .B(_04818_),
    .Y(_04823_));
 sky130_fd_sc_hd__a211o_4 _09848_ (.A1(_04676_),
    .A2(_04822_),
    .B1(_04817_),
    .C1(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__inv_2 _09849_ (.A(_04824_),
    .Y(_01513_));
 sky130_fd_sc_hd__nor2_4 _09850_ (.A(\CPU_Dmem_value_a5[1][26] ),
    .B(_04818_),
    .Y(_04825_));
 sky130_fd_sc_hd__a211o_4 _09851_ (.A1(_04680_),
    .A2(_04822_),
    .B1(_04817_),
    .C1(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__inv_2 _09852_ (.A(_04826_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_4 _09853_ (.A(\CPU_Dmem_value_a5[1][25] ),
    .B(_04818_),
    .Y(_04827_));
 sky130_fd_sc_hd__a211o_4 _09854_ (.A1(_04686_),
    .A2(_04822_),
    .B1(_04817_),
    .C1(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__inv_2 _09855_ (.A(_04828_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_4 _09856_ (.A(\CPU_Dmem_value_a5[1][24] ),
    .B(_04818_),
    .Y(_04829_));
 sky130_fd_sc_hd__a211o_4 _09857_ (.A1(_04690_),
    .A2(_04822_),
    .B1(_04817_),
    .C1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__inv_2 _09858_ (.A(_04830_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_4 _09859_ (.A(\CPU_Dmem_value_a5[1][23] ),
    .B(_04818_),
    .Y(_04831_));
 sky130_fd_sc_hd__a211o_4 _09860_ (.A1(_04695_),
    .A2(_04822_),
    .B1(_04817_),
    .C1(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__inv_2 _09861_ (.A(_04832_),
    .Y(_01509_));
 sky130_fd_sc_hd__buf_2 _09862_ (.A(_04789_),
    .X(_04833_));
 sky130_fd_sc_hd__buf_2 _09863_ (.A(_04808_),
    .X(_04834_));
 sky130_fd_sc_hd__nor2_4 _09864_ (.A(\CPU_Dmem_value_a5[1][22] ),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__a211o_4 _09865_ (.A1(_04699_),
    .A2(_04822_),
    .B1(_04833_),
    .C1(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__inv_2 _09866_ (.A(_04836_),
    .Y(_01508_));
 sky130_fd_sc_hd__buf_2 _09867_ (.A(_04821_),
    .X(_04837_));
 sky130_fd_sc_hd__nor2_4 _09868_ (.A(\CPU_Dmem_value_a5[1][21] ),
    .B(_04834_),
    .Y(_04838_));
 sky130_fd_sc_hd__a211o_4 _09869_ (.A1(_04703_),
    .A2(_04837_),
    .B1(_04833_),
    .C1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__inv_2 _09870_ (.A(_04839_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_4 _09871_ (.A(\CPU_Dmem_value_a5[1][20] ),
    .B(_04834_),
    .Y(_04840_));
 sky130_fd_sc_hd__a211o_4 _09872_ (.A1(_04707_),
    .A2(_04837_),
    .B1(_04833_),
    .C1(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__inv_2 _09873_ (.A(_04841_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_4 _09874_ (.A(\CPU_Dmem_value_a5[1][19] ),
    .B(_04834_),
    .Y(_04842_));
 sky130_fd_sc_hd__a211o_4 _09875_ (.A1(_04713_),
    .A2(_04837_),
    .B1(_04833_),
    .C1(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__inv_2 _09876_ (.A(_04843_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_4 _09877_ (.A(\CPU_Dmem_value_a5[1][18] ),
    .B(_04834_),
    .Y(_04844_));
 sky130_fd_sc_hd__a211o_4 _09878_ (.A1(_04717_),
    .A2(_04837_),
    .B1(_04833_),
    .C1(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__inv_2 _09879_ (.A(_04845_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_4 _09880_ (.A(\CPU_Dmem_value_a5[1][17] ),
    .B(_04834_),
    .Y(_04846_));
 sky130_fd_sc_hd__a211o_4 _09881_ (.A1(_04722_),
    .A2(_04837_),
    .B1(_04833_),
    .C1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__inv_2 _09882_ (.A(_04847_),
    .Y(_01503_));
 sky130_fd_sc_hd__buf_2 _09883_ (.A(_04789_),
    .X(_04848_));
 sky130_fd_sc_hd__buf_2 _09884_ (.A(_04807_),
    .X(_04849_));
 sky130_fd_sc_hd__nor2_4 _09885_ (.A(\CPU_Dmem_value_a5[1][16] ),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__a211o_4 _09886_ (.A1(_04726_),
    .A2(_04837_),
    .B1(_04848_),
    .C1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__inv_2 _09887_ (.A(_04851_),
    .Y(_01502_));
 sky130_fd_sc_hd__buf_2 _09888_ (.A(_04808_),
    .X(_04852_));
 sky130_fd_sc_hd__nor2_4 _09889_ (.A(\CPU_Dmem_value_a5[1][15] ),
    .B(_04849_),
    .Y(_04853_));
 sky130_fd_sc_hd__a211o_4 _09890_ (.A1(_04730_),
    .A2(_04852_),
    .B1(_04848_),
    .C1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__inv_2 _09891_ (.A(_04854_),
    .Y(_01501_));
 sky130_fd_sc_hd__nor2_4 _09892_ (.A(\CPU_Dmem_value_a5[1][14] ),
    .B(_04849_),
    .Y(_04855_));
 sky130_fd_sc_hd__a211o_4 _09893_ (.A1(_04734_),
    .A2(_04852_),
    .B1(_04848_),
    .C1(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__inv_2 _09894_ (.A(_04856_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_4 _09895_ (.A(\CPU_Dmem_value_a5[1][13] ),
    .B(_04849_),
    .Y(_04857_));
 sky130_fd_sc_hd__a211o_4 _09896_ (.A1(_04740_),
    .A2(_04852_),
    .B1(_04848_),
    .C1(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__inv_2 _09897_ (.A(_04858_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_4 _09898_ (.A(\CPU_Dmem_value_a5[1][12] ),
    .B(_04849_),
    .Y(_04859_));
 sky130_fd_sc_hd__a211o_4 _09899_ (.A1(_04744_),
    .A2(_04852_),
    .B1(_04848_),
    .C1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__inv_2 _09900_ (.A(_04860_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_4 _09901_ (.A(\CPU_Dmem_value_a5[1][11] ),
    .B(_04849_),
    .Y(_04861_));
 sky130_fd_sc_hd__a211o_4 _09902_ (.A1(_04749_),
    .A2(_04852_),
    .B1(_04848_),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__inv_2 _09903_ (.A(_04862_),
    .Y(_01497_));
 sky130_fd_sc_hd__buf_2 _09904_ (.A(_04789_),
    .X(_04863_));
 sky130_fd_sc_hd__buf_2 _09905_ (.A(_04807_),
    .X(_04864_));
 sky130_fd_sc_hd__nor2_4 _09906_ (.A(\CPU_Dmem_value_a5[1][10] ),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__a211o_4 _09907_ (.A1(_04753_),
    .A2(_04852_),
    .B1(_04863_),
    .C1(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__inv_2 _09908_ (.A(_04866_),
    .Y(_01496_));
 sky130_fd_sc_hd__buf_2 _09909_ (.A(_04808_),
    .X(_04867_));
 sky130_fd_sc_hd__nor2_4 _09910_ (.A(\CPU_Dmem_value_a5[1][9] ),
    .B(_04864_),
    .Y(_04868_));
 sky130_fd_sc_hd__a211o_4 _09911_ (.A1(_04757_),
    .A2(_04867_),
    .B1(_04863_),
    .C1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__inv_2 _09912_ (.A(_04869_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_4 _09913_ (.A(\CPU_Dmem_value_a5[1][8] ),
    .B(_04864_),
    .Y(_04870_));
 sky130_fd_sc_hd__a211o_4 _09914_ (.A1(_04761_),
    .A2(_04867_),
    .B1(_04863_),
    .C1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__inv_2 _09915_ (.A(_04871_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_4 _09916_ (.A(\CPU_Dmem_value_a5[1][7] ),
    .B(_04864_),
    .Y(_04872_));
 sky130_fd_sc_hd__a211o_4 _09917_ (.A1(_04767_),
    .A2(_04867_),
    .B1(_04863_),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__inv_2 _09918_ (.A(_04873_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_4 _09919_ (.A(\CPU_Dmem_value_a5[1][6] ),
    .B(_04864_),
    .Y(_04874_));
 sky130_fd_sc_hd__a211o_4 _09920_ (.A1(_04771_),
    .A2(_04867_),
    .B1(_04863_),
    .C1(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__inv_2 _09921_ (.A(_04875_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_4 _09922_ (.A(\CPU_Dmem_value_a5[1][5] ),
    .B(_04864_),
    .Y(_04876_));
 sky130_fd_sc_hd__a211o_4 _09923_ (.A1(_04776_),
    .A2(_04867_),
    .B1(_04863_),
    .C1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__inv_2 _09924_ (.A(_04877_),
    .Y(_01491_));
 sky130_fd_sc_hd__buf_2 _09925_ (.A(_04789_),
    .X(_04878_));
 sky130_fd_sc_hd__nor2_4 _09926_ (.A(\CPU_Dmem_value_a5[1][4] ),
    .B(_04821_),
    .Y(_04879_));
 sky130_fd_sc_hd__a211o_4 _09927_ (.A1(_04780_),
    .A2(_04867_),
    .B1(_04878_),
    .C1(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__inv_2 _09928_ (.A(_04880_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_4 _09929_ (.A(\CPU_Dmem_value_a5[1][3] ),
    .B(_04821_),
    .Y(_04881_));
 sky130_fd_sc_hd__a211o_4 _09930_ (.A1(_04784_),
    .A2(_04810_),
    .B1(_04878_),
    .C1(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__inv_2 _09931_ (.A(_04882_),
    .Y(_01489_));
 sky130_fd_sc_hd__nor2_4 _09932_ (.A(\CPU_Dmem_value_a5[1][2] ),
    .B(_04821_),
    .Y(_04883_));
 sky130_fd_sc_hd__a211o_4 _09933_ (.A1(_04788_),
    .A2(_04810_),
    .B1(_04878_),
    .C1(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__inv_2 _09934_ (.A(_04884_),
    .Y(_01488_));
 sky130_fd_sc_hd__nor2_4 _09935_ (.A(\CPU_Dmem_value_a5[1][1] ),
    .B(_04821_),
    .Y(_04885_));
 sky130_fd_sc_hd__a211o_4 _09936_ (.A1(_04794_),
    .A2(_04810_),
    .B1(_04878_),
    .C1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__inv_2 _09937_ (.A(_04886_),
    .Y(_01487_));
 sky130_fd_sc_hd__buf_2 _09938_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .X(_04887_));
 sky130_fd_sc_hd__buf_2 _09939_ (.A(_04660_),
    .X(_04888_));
 sky130_fd_sc_hd__buf_2 _09940_ (.A(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__inv_2 _09941_ (.A(\CPU_Dmem_value_a5[1][0] ),
    .Y(_04890_));
 sky130_fd_sc_hd__nor2_4 _09942_ (.A(_04890_),
    .B(_04809_),
    .Y(_04891_));
 sky130_fd_sc_hd__a211o_4 _09943_ (.A1(_04887_),
    .A2(_04809_),
    .B1(_04889_),
    .C1(_04891_),
    .X(_01486_));
 sky130_fd_sc_hd__inv_2 _09944_ (.A(\CPU_dmem_addr_a4[1] ),
    .Y(_04892_));
 sky130_fd_sc_hd__buf_2 _09945_ (.A(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__or4_4 _09946_ (.A(_04652_),
    .B(_04653_),
    .C(_04893_),
    .D(_04651_),
    .X(_04894_));
 sky130_fd_sc_hd__buf_2 _09947_ (.A(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__nor2_4 _09948_ (.A(_04649_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__buf_2 _09949_ (.A(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__buf_2 _09950_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__buf_2 _09951_ (.A(_04897_),
    .X(_04899_));
 sky130_fd_sc_hd__nor2_4 _09952_ (.A(\CPU_Dmem_value_a5[2][31] ),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__a211o_4 _09953_ (.A1(_04802_),
    .A2(_04898_),
    .B1(_04878_),
    .C1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__inv_2 _09954_ (.A(_04901_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_4 _09955_ (.A(\CPU_Dmem_value_a5[2][30] ),
    .B(_04899_),
    .Y(_04902_));
 sky130_fd_sc_hd__a211o_4 _09956_ (.A1(_04647_),
    .A2(_04898_),
    .B1(_04878_),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__inv_2 _09957_ (.A(_04903_),
    .Y(_01484_));
 sky130_fd_sc_hd__buf_2 _09958_ (.A(CPU_reset_a4),
    .X(_04904_));
 sky130_fd_sc_hd__buf_2 _09959_ (.A(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__buf_2 _09960_ (.A(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__nor2_4 _09961_ (.A(\CPU_Dmem_value_a5[2][29] ),
    .B(_04899_),
    .Y(_04907_));
 sky130_fd_sc_hd__a211o_4 _09962_ (.A1(_04668_),
    .A2(_04898_),
    .B1(_04906_),
    .C1(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__inv_2 _09963_ (.A(_04908_),
    .Y(_01483_));
 sky130_fd_sc_hd__buf_2 _09964_ (.A(_04897_),
    .X(_04909_));
 sky130_fd_sc_hd__nor2_4 _09965_ (.A(\CPU_Dmem_value_a5[2][28] ),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__a211o_4 _09966_ (.A1(_04672_),
    .A2(_04898_),
    .B1(_04906_),
    .C1(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__inv_2 _09967_ (.A(_04911_),
    .Y(_01482_));
 sky130_fd_sc_hd__buf_2 _09968_ (.A(_04896_),
    .X(_04912_));
 sky130_fd_sc_hd__buf_2 _09969_ (.A(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__nor2_4 _09970_ (.A(\CPU_Dmem_value_a5[2][27] ),
    .B(_04909_),
    .Y(_04914_));
 sky130_fd_sc_hd__a211o_4 _09971_ (.A1(_04676_),
    .A2(_04913_),
    .B1(_04906_),
    .C1(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__inv_2 _09972_ (.A(_04915_),
    .Y(_01481_));
 sky130_fd_sc_hd__nor2_4 _09973_ (.A(\CPU_Dmem_value_a5[2][26] ),
    .B(_04909_),
    .Y(_04916_));
 sky130_fd_sc_hd__a211o_4 _09974_ (.A1(_04680_),
    .A2(_04913_),
    .B1(_04906_),
    .C1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__inv_2 _09975_ (.A(_04917_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_4 _09976_ (.A(\CPU_Dmem_value_a5[2][25] ),
    .B(_04909_),
    .Y(_04918_));
 sky130_fd_sc_hd__a211o_4 _09977_ (.A1(_04686_),
    .A2(_04913_),
    .B1(_04906_),
    .C1(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__inv_2 _09978_ (.A(_04919_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_4 _09979_ (.A(\CPU_Dmem_value_a5[2][24] ),
    .B(_04909_),
    .Y(_04920_));
 sky130_fd_sc_hd__a211o_4 _09980_ (.A1(_04690_),
    .A2(_04913_),
    .B1(_04906_),
    .C1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__inv_2 _09981_ (.A(_04921_),
    .Y(_01478_));
 sky130_fd_sc_hd__buf_2 _09982_ (.A(_04905_),
    .X(_04922_));
 sky130_fd_sc_hd__nor2_4 _09983_ (.A(\CPU_Dmem_value_a5[2][23] ),
    .B(_04909_),
    .Y(_04923_));
 sky130_fd_sc_hd__a211o_4 _09984_ (.A1(_04695_),
    .A2(_04913_),
    .B1(_04922_),
    .C1(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__inv_2 _09985_ (.A(_04924_),
    .Y(_01477_));
 sky130_fd_sc_hd__buf_2 _09986_ (.A(_04897_),
    .X(_04925_));
 sky130_fd_sc_hd__nor2_4 _09987_ (.A(\CPU_Dmem_value_a5[2][22] ),
    .B(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__a211o_4 _09988_ (.A1(_04699_),
    .A2(_04913_),
    .B1(_04922_),
    .C1(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__inv_2 _09989_ (.A(_04927_),
    .Y(_01476_));
 sky130_fd_sc_hd__buf_2 _09990_ (.A(_04912_),
    .X(_04928_));
 sky130_fd_sc_hd__nor2_4 _09991_ (.A(\CPU_Dmem_value_a5[2][21] ),
    .B(_04925_),
    .Y(_04929_));
 sky130_fd_sc_hd__a211o_4 _09992_ (.A1(_04703_),
    .A2(_04928_),
    .B1(_04922_),
    .C1(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__inv_2 _09993_ (.A(_04930_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_4 _09994_ (.A(\CPU_Dmem_value_a5[2][20] ),
    .B(_04925_),
    .Y(_04931_));
 sky130_fd_sc_hd__a211o_4 _09995_ (.A1(_04707_),
    .A2(_04928_),
    .B1(_04922_),
    .C1(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__inv_2 _09996_ (.A(_04932_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_4 _09997_ (.A(\CPU_Dmem_value_a5[2][19] ),
    .B(_04925_),
    .Y(_04933_));
 sky130_fd_sc_hd__a211o_4 _09998_ (.A1(_04713_),
    .A2(_04928_),
    .B1(_04922_),
    .C1(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__inv_2 _09999_ (.A(_04934_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_4 _10000_ (.A(\CPU_Dmem_value_a5[2][18] ),
    .B(_04925_),
    .Y(_04935_));
 sky130_fd_sc_hd__a211o_4 _10001_ (.A1(_04717_),
    .A2(_04928_),
    .B1(_04922_),
    .C1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__inv_2 _10002_ (.A(_04936_),
    .Y(_01472_));
 sky130_fd_sc_hd__buf_2 _10003_ (.A(_04905_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_4 _10004_ (.A(\CPU_Dmem_value_a5[2][17] ),
    .B(_04925_),
    .Y(_04938_));
 sky130_fd_sc_hd__a211o_4 _10005_ (.A1(_04722_),
    .A2(_04928_),
    .B1(_04937_),
    .C1(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__inv_2 _10006_ (.A(_04939_),
    .Y(_01471_));
 sky130_fd_sc_hd__buf_2 _10007_ (.A(_04896_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_4 _10008_ (.A(\CPU_Dmem_value_a5[2][16] ),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__a211o_4 _10009_ (.A1(_04726_),
    .A2(_04928_),
    .B1(_04937_),
    .C1(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__inv_2 _10010_ (.A(_04942_),
    .Y(_01470_));
 sky130_fd_sc_hd__buf_2 _10011_ (.A(_04897_),
    .X(_04943_));
 sky130_fd_sc_hd__nor2_4 _10012_ (.A(\CPU_Dmem_value_a5[2][15] ),
    .B(_04940_),
    .Y(_04944_));
 sky130_fd_sc_hd__a211o_4 _10013_ (.A1(_04730_),
    .A2(_04943_),
    .B1(_04937_),
    .C1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__inv_2 _10014_ (.A(_04945_),
    .Y(_01469_));
 sky130_fd_sc_hd__nor2_4 _10015_ (.A(\CPU_Dmem_value_a5[2][14] ),
    .B(_04940_),
    .Y(_04946_));
 sky130_fd_sc_hd__a211o_4 _10016_ (.A1(_04734_),
    .A2(_04943_),
    .B1(_04937_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__inv_2 _10017_ (.A(_04947_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_4 _10018_ (.A(\CPU_Dmem_value_a5[2][13] ),
    .B(_04940_),
    .Y(_04948_));
 sky130_fd_sc_hd__a211o_4 _10019_ (.A1(_04740_),
    .A2(_04943_),
    .B1(_04937_),
    .C1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__inv_2 _10020_ (.A(_04949_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_4 _10021_ (.A(\CPU_Dmem_value_a5[2][12] ),
    .B(_04940_),
    .Y(_04950_));
 sky130_fd_sc_hd__a211o_4 _10022_ (.A1(_04744_),
    .A2(_04943_),
    .B1(_04937_),
    .C1(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__inv_2 _10023_ (.A(_04951_),
    .Y(_01466_));
 sky130_fd_sc_hd__buf_2 _10024_ (.A(_04905_),
    .X(_04952_));
 sky130_fd_sc_hd__nor2_4 _10025_ (.A(\CPU_Dmem_value_a5[2][11] ),
    .B(_04940_),
    .Y(_04953_));
 sky130_fd_sc_hd__a211o_4 _10026_ (.A1(_04749_),
    .A2(_04943_),
    .B1(_04952_),
    .C1(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__inv_2 _10027_ (.A(_04954_),
    .Y(_01465_));
 sky130_fd_sc_hd__buf_2 _10028_ (.A(_04896_),
    .X(_04955_));
 sky130_fd_sc_hd__nor2_4 _10029_ (.A(\CPU_Dmem_value_a5[2][10] ),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__a211o_4 _10030_ (.A1(_04753_),
    .A2(_04943_),
    .B1(_04952_),
    .C1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__inv_2 _10031_ (.A(_04957_),
    .Y(_01464_));
 sky130_fd_sc_hd__buf_2 _10032_ (.A(_04897_),
    .X(_04958_));
 sky130_fd_sc_hd__nor2_4 _10033_ (.A(\CPU_Dmem_value_a5[2][9] ),
    .B(_04955_),
    .Y(_04959_));
 sky130_fd_sc_hd__a211o_4 _10034_ (.A1(_04757_),
    .A2(_04958_),
    .B1(_04952_),
    .C1(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__inv_2 _10035_ (.A(_04960_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_4 _10036_ (.A(\CPU_Dmem_value_a5[2][8] ),
    .B(_04955_),
    .Y(_04961_));
 sky130_fd_sc_hd__a211o_4 _10037_ (.A1(_04761_),
    .A2(_04958_),
    .B1(_04952_),
    .C1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__inv_2 _10038_ (.A(_04962_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_4 _10039_ (.A(\CPU_Dmem_value_a5[2][7] ),
    .B(_04955_),
    .Y(_04963_));
 sky130_fd_sc_hd__a211o_4 _10040_ (.A1(_04767_),
    .A2(_04958_),
    .B1(_04952_),
    .C1(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__inv_2 _10041_ (.A(_04964_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_4 _10042_ (.A(\CPU_Dmem_value_a5[2][6] ),
    .B(_04955_),
    .Y(_04965_));
 sky130_fd_sc_hd__a211o_4 _10043_ (.A1(_04771_),
    .A2(_04958_),
    .B1(_04952_),
    .C1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__inv_2 _10044_ (.A(_04966_),
    .Y(_01460_));
 sky130_fd_sc_hd__buf_2 _10045_ (.A(_04905_),
    .X(_04967_));
 sky130_fd_sc_hd__nor2_4 _10046_ (.A(\CPU_Dmem_value_a5[2][5] ),
    .B(_04955_),
    .Y(_04968_));
 sky130_fd_sc_hd__a211o_4 _10047_ (.A1(_04776_),
    .A2(_04958_),
    .B1(_04967_),
    .C1(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__inv_2 _10048_ (.A(_04969_),
    .Y(_01459_));
 sky130_fd_sc_hd__nor2_4 _10049_ (.A(\CPU_Dmem_value_a5[2][4] ),
    .B(_04912_),
    .Y(_04970_));
 sky130_fd_sc_hd__a211o_4 _10050_ (.A1(_04780_),
    .A2(_04958_),
    .B1(_04967_),
    .C1(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__inv_2 _10051_ (.A(_04971_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_4 _10052_ (.A(\CPU_Dmem_value_a5[2][3] ),
    .B(_04912_),
    .Y(_04972_));
 sky130_fd_sc_hd__a211o_4 _10053_ (.A1(_04784_),
    .A2(_04899_),
    .B1(_04967_),
    .C1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__inv_2 _10054_ (.A(_04973_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_4 _10055_ (.A(\CPU_Dmem_value_a5[2][2] ),
    .B(_04912_),
    .Y(_04974_));
 sky130_fd_sc_hd__a211o_4 _10056_ (.A1(_04788_),
    .A2(_04899_),
    .B1(_04967_),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__inv_2 _10057_ (.A(_04975_),
    .Y(_01456_));
 sky130_fd_sc_hd__buf_2 _10058_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .X(_04976_));
 sky130_fd_sc_hd__inv_2 _10059_ (.A(\CPU_Dmem_value_a5[2][1] ),
    .Y(_04977_));
 sky130_fd_sc_hd__nor2_4 _10060_ (.A(_04977_),
    .B(_04898_),
    .Y(_04978_));
 sky130_fd_sc_hd__a211o_4 _10061_ (.A1(_04976_),
    .A2(_04898_),
    .B1(_04889_),
    .C1(_04978_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2_4 _10062_ (.A(\CPU_Dmem_value_a5[2][0] ),
    .B(_04912_),
    .Y(_04979_));
 sky130_fd_sc_hd__a211o_4 _10063_ (.A1(_04798_),
    .A2(_04899_),
    .B1(_04967_),
    .C1(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__inv_2 _10064_ (.A(_04980_),
    .Y(_01454_));
 sky130_fd_sc_hd__or4_4 _10065_ (.A(_04652_),
    .B(_04653_),
    .C(_04893_),
    .D(_04804_),
    .X(_04981_));
 sky130_fd_sc_hd__buf_2 _10066_ (.A(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__nor2_4 _10067_ (.A(_04649_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__buf_2 _10068_ (.A(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__buf_2 _10069_ (.A(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__buf_2 _10070_ (.A(_04984_),
    .X(_04986_));
 sky130_fd_sc_hd__nor2_4 _10071_ (.A(\CPU_Dmem_value_a5[3][31] ),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__a211o_4 _10072_ (.A1(_04802_),
    .A2(_04985_),
    .B1(_04967_),
    .C1(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__inv_2 _10073_ (.A(_04988_),
    .Y(_01453_));
 sky130_fd_sc_hd__buf_2 _10074_ (.A(_04905_),
    .X(_04989_));
 sky130_fd_sc_hd__nor2_4 _10075_ (.A(\CPU_Dmem_value_a5[3][30] ),
    .B(_04986_),
    .Y(_04990_));
 sky130_fd_sc_hd__a211o_4 _10076_ (.A1(_04647_),
    .A2(_04985_),
    .B1(_04989_),
    .C1(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__inv_2 _10077_ (.A(_04991_),
    .Y(_01452_));
 sky130_fd_sc_hd__buf_2 _10078_ (.A(_04983_),
    .X(_04992_));
 sky130_fd_sc_hd__buf_2 _10079_ (.A(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__buf_2 _10080_ (.A(_04984_),
    .X(_04994_));
 sky130_fd_sc_hd__nor2_4 _10081_ (.A(\CPU_Dmem_value_a5[3][29] ),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__a211o_4 _10082_ (.A1(_04668_),
    .A2(_04993_),
    .B1(_04989_),
    .C1(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__inv_2 _10083_ (.A(_04996_),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_4 _10084_ (.A(\CPU_Dmem_value_a5[3][28] ),
    .B(_04994_),
    .Y(_04997_));
 sky130_fd_sc_hd__a211o_4 _10085_ (.A1(_04672_),
    .A2(_04993_),
    .B1(_04989_),
    .C1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__inv_2 _10086_ (.A(_04998_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_4 _10087_ (.A(\CPU_Dmem_value_a5[3][27] ),
    .B(_04994_),
    .Y(_04999_));
 sky130_fd_sc_hd__a211o_4 _10088_ (.A1(_04676_),
    .A2(_04993_),
    .B1(_04989_),
    .C1(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__inv_2 _10089_ (.A(_05000_),
    .Y(_01449_));
 sky130_fd_sc_hd__nor2_4 _10090_ (.A(\CPU_Dmem_value_a5[3][26] ),
    .B(_04994_),
    .Y(_05001_));
 sky130_fd_sc_hd__a211o_4 _10091_ (.A1(_04680_),
    .A2(_04993_),
    .B1(_04989_),
    .C1(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__inv_2 _10092_ (.A(_05002_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_4 _10093_ (.A(\CPU_Dmem_value_a5[3][25] ),
    .B(_04994_),
    .Y(_05003_));
 sky130_fd_sc_hd__a211o_4 _10094_ (.A1(_04686_),
    .A2(_04993_),
    .B1(_04989_),
    .C1(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__inv_2 _10095_ (.A(_05004_),
    .Y(_01447_));
 sky130_fd_sc_hd__buf_2 _10096_ (.A(_04904_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_2 _10097_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__nor2_4 _10098_ (.A(\CPU_Dmem_value_a5[3][24] ),
    .B(_04994_),
    .Y(_05007_));
 sky130_fd_sc_hd__a211o_4 _10099_ (.A1(_04690_),
    .A2(_04993_),
    .B1(_05006_),
    .C1(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__inv_2 _10100_ (.A(_05008_),
    .Y(_01446_));
 sky130_fd_sc_hd__buf_2 _10101_ (.A(_04992_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_2 _10102_ (.A(_04984_),
    .X(_05010_));
 sky130_fd_sc_hd__nor2_4 _10103_ (.A(\CPU_Dmem_value_a5[3][23] ),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__a211o_4 _10104_ (.A1(_04695_),
    .A2(_05009_),
    .B1(_05006_),
    .C1(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_05012_),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_4 _10106_ (.A(\CPU_Dmem_value_a5[3][22] ),
    .B(_05010_),
    .Y(_05013_));
 sky130_fd_sc_hd__a211o_4 _10107_ (.A1(_04699_),
    .A2(_05009_),
    .B1(_05006_),
    .C1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__inv_2 _10108_ (.A(_05014_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_4 _10109_ (.A(\CPU_Dmem_value_a5[3][21] ),
    .B(_05010_),
    .Y(_05015_));
 sky130_fd_sc_hd__a211o_4 _10110_ (.A1(_04703_),
    .A2(_05009_),
    .B1(_05006_),
    .C1(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__inv_2 _10111_ (.A(_05016_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_4 _10112_ (.A(\CPU_Dmem_value_a5[3][20] ),
    .B(_05010_),
    .Y(_05017_));
 sky130_fd_sc_hd__a211o_4 _10113_ (.A1(_04707_),
    .A2(_05009_),
    .B1(_05006_),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__inv_2 _10114_ (.A(_05018_),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_4 _10115_ (.A(\CPU_Dmem_value_a5[3][19] ),
    .B(_05010_),
    .Y(_05019_));
 sky130_fd_sc_hd__a211o_4 _10116_ (.A1(_04713_),
    .A2(_05009_),
    .B1(_05006_),
    .C1(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__inv_2 _10117_ (.A(_05020_),
    .Y(_01441_));
 sky130_fd_sc_hd__buf_2 _10118_ (.A(_05005_),
    .X(_05021_));
 sky130_fd_sc_hd__nor2_4 _10119_ (.A(\CPU_Dmem_value_a5[3][18] ),
    .B(_05010_),
    .Y(_05022_));
 sky130_fd_sc_hd__a211o_4 _10120_ (.A1(_04717_),
    .A2(_05009_),
    .B1(_05021_),
    .C1(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__inv_2 _10121_ (.A(_05023_),
    .Y(_01440_));
 sky130_fd_sc_hd__buf_2 _10122_ (.A(_04984_),
    .X(_05024_));
 sky130_fd_sc_hd__buf_2 _10123_ (.A(_04983_),
    .X(_05025_));
 sky130_fd_sc_hd__nor2_4 _10124_ (.A(\CPU_Dmem_value_a5[3][17] ),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__a211o_4 _10125_ (.A1(_04722_),
    .A2(_05024_),
    .B1(_05021_),
    .C1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__inv_2 _10126_ (.A(_05027_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_4 _10127_ (.A(\CPU_Dmem_value_a5[3][16] ),
    .B(_05025_),
    .Y(_05028_));
 sky130_fd_sc_hd__a211o_4 _10128_ (.A1(_04726_),
    .A2(_05024_),
    .B1(_05021_),
    .C1(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__inv_2 _10129_ (.A(_05029_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_4 _10130_ (.A(\CPU_Dmem_value_a5[3][15] ),
    .B(_05025_),
    .Y(_05030_));
 sky130_fd_sc_hd__a211o_4 _10131_ (.A1(_04730_),
    .A2(_05024_),
    .B1(_05021_),
    .C1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__inv_2 _10132_ (.A(_05031_),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_4 _10133_ (.A(\CPU_Dmem_value_a5[3][14] ),
    .B(_05025_),
    .Y(_05032_));
 sky130_fd_sc_hd__a211o_4 _10134_ (.A1(_04734_),
    .A2(_05024_),
    .B1(_05021_),
    .C1(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__inv_2 _10135_ (.A(_05033_),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_4 _10136_ (.A(\CPU_Dmem_value_a5[3][13] ),
    .B(_05025_),
    .Y(_05034_));
 sky130_fd_sc_hd__a211o_4 _10137_ (.A1(_04740_),
    .A2(_05024_),
    .B1(_05021_),
    .C1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__inv_2 _10138_ (.A(_05035_),
    .Y(_01435_));
 sky130_fd_sc_hd__buf_2 _10139_ (.A(_05005_),
    .X(_05036_));
 sky130_fd_sc_hd__nor2_4 _10140_ (.A(\CPU_Dmem_value_a5[3][12] ),
    .B(_05025_),
    .Y(_05037_));
 sky130_fd_sc_hd__a211o_4 _10141_ (.A1(_04744_),
    .A2(_05024_),
    .B1(_05036_),
    .C1(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__inv_2 _10142_ (.A(_05038_),
    .Y(_01434_));
 sky130_fd_sc_hd__buf_2 _10143_ (.A(_04984_),
    .X(_05039_));
 sky130_fd_sc_hd__buf_2 _10144_ (.A(_04983_),
    .X(_05040_));
 sky130_fd_sc_hd__nor2_4 _10145_ (.A(\CPU_Dmem_value_a5[3][11] ),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a211o_4 _10146_ (.A1(_04749_),
    .A2(_05039_),
    .B1(_05036_),
    .C1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_05042_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_4 _10148_ (.A(\CPU_Dmem_value_a5[3][10] ),
    .B(_05040_),
    .Y(_05043_));
 sky130_fd_sc_hd__a211o_4 _10149_ (.A1(_04753_),
    .A2(_05039_),
    .B1(_05036_),
    .C1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__inv_2 _10150_ (.A(_05044_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_4 _10151_ (.A(\CPU_Dmem_value_a5[3][9] ),
    .B(_05040_),
    .Y(_05045_));
 sky130_fd_sc_hd__a211o_4 _10152_ (.A1(_04757_),
    .A2(_05039_),
    .B1(_05036_),
    .C1(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__inv_2 _10153_ (.A(_05046_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_4 _10154_ (.A(\CPU_Dmem_value_a5[3][8] ),
    .B(_05040_),
    .Y(_05047_));
 sky130_fd_sc_hd__a211o_4 _10155_ (.A1(_04761_),
    .A2(_05039_),
    .B1(_05036_),
    .C1(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__inv_2 _10156_ (.A(_05048_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_4 _10157_ (.A(\CPU_Dmem_value_a5[3][7] ),
    .B(_05040_),
    .Y(_05049_));
 sky130_fd_sc_hd__a211o_4 _10158_ (.A1(_04767_),
    .A2(_05039_),
    .B1(_05036_),
    .C1(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__inv_2 _10159_ (.A(_05050_),
    .Y(_01429_));
 sky130_fd_sc_hd__buf_2 _10160_ (.A(_05005_),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_4 _10161_ (.A(\CPU_Dmem_value_a5[3][6] ),
    .B(_05040_),
    .Y(_05052_));
 sky130_fd_sc_hd__a211o_4 _10162_ (.A1(_04771_),
    .A2(_05039_),
    .B1(_05051_),
    .C1(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__inv_2 _10163_ (.A(_05053_),
    .Y(_01428_));
 sky130_fd_sc_hd__nor2_4 _10164_ (.A(\CPU_Dmem_value_a5[3][5] ),
    .B(_04992_),
    .Y(_05054_));
 sky130_fd_sc_hd__a211o_4 _10165_ (.A1(_04776_),
    .A2(_04986_),
    .B1(_05051_),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__inv_2 _10166_ (.A(_05055_),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_4 _10167_ (.A(\CPU_Dmem_value_a5[3][4] ),
    .B(_04992_),
    .Y(_05056_));
 sky130_fd_sc_hd__a211o_4 _10168_ (.A1(_04780_),
    .A2(_04986_),
    .B1(_05051_),
    .C1(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__inv_2 _10169_ (.A(_05057_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_4 _10170_ (.A(\CPU_Dmem_value_a5[3][3] ),
    .B(_04992_),
    .Y(_05058_));
 sky130_fd_sc_hd__a211o_4 _10171_ (.A1(_04784_),
    .A2(_04986_),
    .B1(_05051_),
    .C1(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__inv_2 _10172_ (.A(_05059_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_4 _10173_ (.A(\CPU_Dmem_value_a5[3][2] ),
    .B(_04992_),
    .Y(_05060_));
 sky130_fd_sc_hd__a211o_4 _10174_ (.A1(_04788_),
    .A2(_04986_),
    .B1(_05051_),
    .C1(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__inv_2 _10175_ (.A(_05061_),
    .Y(_01424_));
 sky130_fd_sc_hd__inv_2 _10176_ (.A(\CPU_Dmem_value_a5[3][1] ),
    .Y(_05062_));
 sky130_fd_sc_hd__nor2_4 _10177_ (.A(_05062_),
    .B(_04985_),
    .Y(_05063_));
 sky130_fd_sc_hd__a211o_4 _10178_ (.A1(_04976_),
    .A2(_04985_),
    .B1(_04889_),
    .C1(_05063_),
    .X(_01423_));
 sky130_fd_sc_hd__inv_2 _10179_ (.A(\CPU_Dmem_value_a5[3][0] ),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_4 _10180_ (.A(_05064_),
    .B(_04985_),
    .Y(_05065_));
 sky130_fd_sc_hd__a211o_4 _10181_ (.A1(_04887_),
    .A2(_04985_),
    .B1(_04889_),
    .C1(_05065_),
    .X(_01422_));
 sky130_fd_sc_hd__inv_2 _10182_ (.A(\CPU_dmem_addr_a4[2] ),
    .Y(_05066_));
 sky130_fd_sc_hd__buf_2 _10183_ (.A(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__or4_4 _10184_ (.A(_04650_),
    .B(_04651_),
    .C(_04652_),
    .D(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__or2_4 _10185_ (.A(_04648_),
    .B(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__inv_2 _10186_ (.A(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__buf_2 _10187_ (.A(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__buf_2 _10188_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__buf_2 _10189_ (.A(_05070_),
    .X(_05073_));
 sky130_fd_sc_hd__buf_2 _10190_ (.A(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__nor2_4 _10191_ (.A(\CPU_Dmem_value_a5[4][31] ),
    .B(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__a211o_4 _10192_ (.A1(_04802_),
    .A2(_05072_),
    .B1(_05051_),
    .C1(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__inv_2 _10193_ (.A(_05076_),
    .Y(_01421_));
 sky130_fd_sc_hd__buf_2 _10194_ (.A(_05005_),
    .X(_05077_));
 sky130_fd_sc_hd__nor2_4 _10195_ (.A(\CPU_Dmem_value_a5[4][30] ),
    .B(_05074_),
    .Y(_05078_));
 sky130_fd_sc_hd__a211o_4 _10196_ (.A1(_04647_),
    .A2(_05072_),
    .B1(_05077_),
    .C1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__inv_2 _10197_ (.A(_05079_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_4 _10198_ (.A(\CPU_Dmem_value_a5[4][29] ),
    .B(_05074_),
    .Y(_05080_));
 sky130_fd_sc_hd__a211o_4 _10199_ (.A1(_04668_),
    .A2(_05072_),
    .B1(_05077_),
    .C1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__inv_2 _10200_ (.A(_05081_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_4 _10201_ (.A(\CPU_Dmem_value_a5[4][28] ),
    .B(_05074_),
    .Y(_05082_));
 sky130_fd_sc_hd__a211o_4 _10202_ (.A1(_04672_),
    .A2(_05072_),
    .B1(_05077_),
    .C1(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__inv_2 _10203_ (.A(_05083_),
    .Y(_01418_));
 sky130_fd_sc_hd__buf_2 _10204_ (.A(_05073_),
    .X(_05084_));
 sky130_fd_sc_hd__nor2_4 _10205_ (.A(\CPU_Dmem_value_a5[4][27] ),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a211o_4 _10206_ (.A1(_04676_),
    .A2(_05072_),
    .B1(_05077_),
    .C1(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__inv_2 _10207_ (.A(_05086_),
    .Y(_01417_));
 sky130_fd_sc_hd__buf_2 _10208_ (.A(_05071_),
    .X(_05087_));
 sky130_fd_sc_hd__nor2_4 _10209_ (.A(\CPU_Dmem_value_a5[4][26] ),
    .B(_05084_),
    .Y(_05088_));
 sky130_fd_sc_hd__a211o_4 _10210_ (.A1(_04680_),
    .A2(_05087_),
    .B1(_05077_),
    .C1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__inv_2 _10211_ (.A(_05089_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_4 _10212_ (.A(\CPU_Dmem_value_a5[4][25] ),
    .B(_05084_),
    .Y(_05090_));
 sky130_fd_sc_hd__a211o_4 _10213_ (.A1(_04686_),
    .A2(_05087_),
    .B1(_05077_),
    .C1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__inv_2 _10214_ (.A(_05091_),
    .Y(_01415_));
 sky130_fd_sc_hd__buf_2 _10215_ (.A(_05005_),
    .X(_05092_));
 sky130_fd_sc_hd__nor2_4 _10216_ (.A(\CPU_Dmem_value_a5[4][24] ),
    .B(_05084_),
    .Y(_05093_));
 sky130_fd_sc_hd__a211o_4 _10217_ (.A1(_04690_),
    .A2(_05087_),
    .B1(_05092_),
    .C1(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__inv_2 _10218_ (.A(_05094_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_4 _10219_ (.A(\CPU_Dmem_value_a5[4][23] ),
    .B(_05084_),
    .Y(_05095_));
 sky130_fd_sc_hd__a211o_4 _10220_ (.A1(_04695_),
    .A2(_05087_),
    .B1(_05092_),
    .C1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__inv_2 _10221_ (.A(_05096_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_4 _10222_ (.A(\CPU_Dmem_value_a5[4][22] ),
    .B(_05084_),
    .Y(_05097_));
 sky130_fd_sc_hd__a211o_4 _10223_ (.A1(_04699_),
    .A2(_05087_),
    .B1(_05092_),
    .C1(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__inv_2 _10224_ (.A(_05098_),
    .Y(_01412_));
 sky130_fd_sc_hd__buf_2 _10225_ (.A(_05073_),
    .X(_05099_));
 sky130_fd_sc_hd__nor2_4 _10226_ (.A(\CPU_Dmem_value_a5[4][21] ),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__a211o_4 _10227_ (.A1(_04703_),
    .A2(_05087_),
    .B1(_05092_),
    .C1(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__inv_2 _10228_ (.A(_05101_),
    .Y(_01411_));
 sky130_fd_sc_hd__buf_2 _10229_ (.A(_05071_),
    .X(_05102_));
 sky130_fd_sc_hd__nor2_4 _10230_ (.A(\CPU_Dmem_value_a5[4][20] ),
    .B(_05099_),
    .Y(_05103_));
 sky130_fd_sc_hd__a211o_4 _10231_ (.A1(_04707_),
    .A2(_05102_),
    .B1(_05092_),
    .C1(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__inv_2 _10232_ (.A(_05104_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_4 _10233_ (.A(\CPU_Dmem_value_a5[4][19] ),
    .B(_05099_),
    .Y(_05105_));
 sky130_fd_sc_hd__a211o_4 _10234_ (.A1(_04713_),
    .A2(_05102_),
    .B1(_05092_),
    .C1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__inv_2 _10235_ (.A(_05106_),
    .Y(_01409_));
 sky130_fd_sc_hd__buf_2 _10236_ (.A(_04904_),
    .X(_05107_));
 sky130_fd_sc_hd__buf_2 _10237_ (.A(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_4 _10238_ (.A(\CPU_Dmem_value_a5[4][18] ),
    .B(_05099_),
    .Y(_05109_));
 sky130_fd_sc_hd__a211o_4 _10239_ (.A1(_04717_),
    .A2(_05102_),
    .B1(_05108_),
    .C1(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__inv_2 _10240_ (.A(_05110_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_4 _10241_ (.A(\CPU_Dmem_value_a5[4][17] ),
    .B(_05099_),
    .Y(_05111_));
 sky130_fd_sc_hd__a211o_4 _10242_ (.A1(_04722_),
    .A2(_05102_),
    .B1(_05108_),
    .C1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__inv_2 _10243_ (.A(_05112_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_4 _10244_ (.A(\CPU_Dmem_value_a5[4][16] ),
    .B(_05099_),
    .Y(_05113_));
 sky130_fd_sc_hd__a211o_4 _10245_ (.A1(_04726_),
    .A2(_05102_),
    .B1(_05108_),
    .C1(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__inv_2 _10246_ (.A(_05114_),
    .Y(_01406_));
 sky130_fd_sc_hd__buf_2 _10247_ (.A(_05073_),
    .X(_05115_));
 sky130_fd_sc_hd__nor2_4 _10248_ (.A(\CPU_Dmem_value_a5[4][15] ),
    .B(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__a211o_4 _10249_ (.A1(_04730_),
    .A2(_05102_),
    .B1(_05108_),
    .C1(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__inv_2 _10250_ (.A(_05117_),
    .Y(_01405_));
 sky130_fd_sc_hd__buf_2 _10251_ (.A(_05071_),
    .X(_05118_));
 sky130_fd_sc_hd__nor2_4 _10252_ (.A(\CPU_Dmem_value_a5[4][14] ),
    .B(_05115_),
    .Y(_05119_));
 sky130_fd_sc_hd__a211o_4 _10253_ (.A1(_04734_),
    .A2(_05118_),
    .B1(_05108_),
    .C1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__inv_2 _10254_ (.A(_05120_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_4 _10255_ (.A(\CPU_Dmem_value_a5[4][13] ),
    .B(_05115_),
    .Y(_05121_));
 sky130_fd_sc_hd__a211o_4 _10256_ (.A1(_04740_),
    .A2(_05118_),
    .B1(_05108_),
    .C1(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__inv_2 _10257_ (.A(_05122_),
    .Y(_01403_));
 sky130_fd_sc_hd__buf_2 _10258_ (.A(_05107_),
    .X(_05123_));
 sky130_fd_sc_hd__nor2_4 _10259_ (.A(\CPU_Dmem_value_a5[4][12] ),
    .B(_05115_),
    .Y(_05124_));
 sky130_fd_sc_hd__a211o_4 _10260_ (.A1(_04744_),
    .A2(_05118_),
    .B1(_05123_),
    .C1(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__inv_2 _10261_ (.A(_05125_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_4 _10262_ (.A(\CPU_Dmem_value_a5[4][11] ),
    .B(_05115_),
    .Y(_05126_));
 sky130_fd_sc_hd__a211o_4 _10263_ (.A1(_04749_),
    .A2(_05118_),
    .B1(_05123_),
    .C1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__inv_2 _10264_ (.A(_05127_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_4 _10265_ (.A(\CPU_Dmem_value_a5[4][10] ),
    .B(_05115_),
    .Y(_05128_));
 sky130_fd_sc_hd__a211o_4 _10266_ (.A1(_04753_),
    .A2(_05118_),
    .B1(_05123_),
    .C1(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__inv_2 _10267_ (.A(_05129_),
    .Y(_01400_));
 sky130_fd_sc_hd__buf_2 _10268_ (.A(_05073_),
    .X(_05130_));
 sky130_fd_sc_hd__nor2_4 _10269_ (.A(\CPU_Dmem_value_a5[4][9] ),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__a211o_4 _10270_ (.A1(_04757_),
    .A2(_05118_),
    .B1(_05123_),
    .C1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__inv_2 _10271_ (.A(_05132_),
    .Y(_01399_));
 sky130_fd_sc_hd__buf_2 _10272_ (.A(_05073_),
    .X(_05133_));
 sky130_fd_sc_hd__nor2_4 _10273_ (.A(\CPU_Dmem_value_a5[4][8] ),
    .B(_05130_),
    .Y(_05134_));
 sky130_fd_sc_hd__a211o_4 _10274_ (.A1(_04761_),
    .A2(_05133_),
    .B1(_05123_),
    .C1(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__inv_2 _10275_ (.A(_05135_),
    .Y(_01398_));
 sky130_fd_sc_hd__nor2_4 _10276_ (.A(\CPU_Dmem_value_a5[4][7] ),
    .B(_05130_),
    .Y(_05136_));
 sky130_fd_sc_hd__a211o_4 _10277_ (.A1(_04767_),
    .A2(_05133_),
    .B1(_05123_),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__inv_2 _10278_ (.A(_05137_),
    .Y(_01397_));
 sky130_fd_sc_hd__buf_2 _10279_ (.A(_05107_),
    .X(_05138_));
 sky130_fd_sc_hd__nor2_4 _10280_ (.A(\CPU_Dmem_value_a5[4][6] ),
    .B(_05130_),
    .Y(_05139_));
 sky130_fd_sc_hd__a211o_4 _10281_ (.A1(_04771_),
    .A2(_05133_),
    .B1(_05138_),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__inv_2 _10282_ (.A(_05140_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_4 _10283_ (.A(\CPU_Dmem_value_a5[4][5] ),
    .B(_05130_),
    .Y(_05141_));
 sky130_fd_sc_hd__a211o_4 _10284_ (.A1(_04776_),
    .A2(_05133_),
    .B1(_05138_),
    .C1(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__inv_2 _10285_ (.A(_05142_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_4 _10286_ (.A(\CPU_Dmem_value_a5[4][4] ),
    .B(_05130_),
    .Y(_05143_));
 sky130_fd_sc_hd__a211o_4 _10287_ (.A1(_04780_),
    .A2(_05133_),
    .B1(_05138_),
    .C1(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__inv_2 _10288_ (.A(_05144_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_4 _10289_ (.A(\CPU_Dmem_value_a5[4][3] ),
    .B(_05071_),
    .Y(_05145_));
 sky130_fd_sc_hd__a211o_4 _10290_ (.A1(_04784_),
    .A2(_05133_),
    .B1(_05138_),
    .C1(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__inv_2 _10291_ (.A(_05146_),
    .Y(_01393_));
 sky130_fd_sc_hd__buf_2 _10292_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .X(_05147_));
 sky130_fd_sc_hd__and2_4 _10293_ (.A(\CPU_Dmem_value_a5[4][2] ),
    .B(_05069_),
    .X(_05148_));
 sky130_fd_sc_hd__a211o_4 _10294_ (.A1(_05147_),
    .A2(_05072_),
    .B1(_04889_),
    .C1(_05148_),
    .X(_01392_));
 sky130_fd_sc_hd__nor2_4 _10295_ (.A(\CPU_Dmem_value_a5[4][1] ),
    .B(_05071_),
    .Y(_05149_));
 sky130_fd_sc_hd__a211o_4 _10296_ (.A1(_04794_),
    .A2(_05074_),
    .B1(_05138_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__inv_2 _10297_ (.A(_05150_),
    .Y(_01391_));
 sky130_fd_sc_hd__inv_2 _10298_ (.A(\CPU_Dmem_value_a5[4][0] ),
    .Y(_05151_));
 sky130_fd_sc_hd__and2_4 _10299_ (.A(_05151_),
    .B(_05069_),
    .X(_05152_));
 sky130_fd_sc_hd__a211o_4 _10300_ (.A1(_04798_),
    .A2(_05074_),
    .B1(_05138_),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__inv_2 _10301_ (.A(_05153_),
    .Y(_01390_));
 sky130_fd_sc_hd__or4_4 _10302_ (.A(_04650_),
    .B(_04804_),
    .C(_04652_),
    .D(_05067_),
    .X(_05154_));
 sky130_fd_sc_hd__or2_4 _10303_ (.A(_04648_),
    .B(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__inv_2 _10304_ (.A(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__buf_2 _10305_ (.A(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__buf_2 _10306_ (.A(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__buf_2 _10307_ (.A(_05107_),
    .X(_05159_));
 sky130_fd_sc_hd__buf_2 _10308_ (.A(_05156_),
    .X(_05160_));
 sky130_fd_sc_hd__buf_2 _10309_ (.A(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_4 _10310_ (.A(\CPU_Dmem_value_a5[5][31] ),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__a211o_4 _10311_ (.A1(_04802_),
    .A2(_05158_),
    .B1(_05159_),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__inv_2 _10312_ (.A(_05163_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_4 _10313_ (.A(\CPU_Dmem_value_a5[5][30] ),
    .B(_05161_),
    .Y(_05164_));
 sky130_fd_sc_hd__a211o_4 _10314_ (.A1(_04647_),
    .A2(_05158_),
    .B1(_05159_),
    .C1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__inv_2 _10315_ (.A(_05165_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_4 _10316_ (.A(\CPU_Dmem_value_a5[5][29] ),
    .B(_05161_),
    .Y(_05166_));
 sky130_fd_sc_hd__a211o_4 _10317_ (.A1(_04668_),
    .A2(_05158_),
    .B1(_05159_),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__inv_2 _10318_ (.A(_05167_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_4 _10319_ (.A(\CPU_Dmem_value_a5[5][28] ),
    .B(_05161_),
    .Y(_05168_));
 sky130_fd_sc_hd__a211o_4 _10320_ (.A1(_04672_),
    .A2(_05158_),
    .B1(_05159_),
    .C1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__inv_2 _10321_ (.A(_05169_),
    .Y(_01386_));
 sky130_fd_sc_hd__buf_2 _10322_ (.A(_05157_),
    .X(_05170_));
 sky130_fd_sc_hd__buf_2 _10323_ (.A(_05160_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_4 _10324_ (.A(\CPU_Dmem_value_a5[5][27] ),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a211o_4 _10325_ (.A1(_04676_),
    .A2(_05170_),
    .B1(_05159_),
    .C1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__inv_2 _10326_ (.A(_05173_),
    .Y(_01385_));
 sky130_fd_sc_hd__nor2_4 _10327_ (.A(\CPU_Dmem_value_a5[5][26] ),
    .B(_05171_),
    .Y(_05174_));
 sky130_fd_sc_hd__a211o_4 _10328_ (.A1(_04680_),
    .A2(_05170_),
    .B1(_05159_),
    .C1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__inv_2 _10329_ (.A(_05175_),
    .Y(_01384_));
 sky130_fd_sc_hd__buf_2 _10330_ (.A(_05107_),
    .X(_05176_));
 sky130_fd_sc_hd__nor2_4 _10331_ (.A(\CPU_Dmem_value_a5[5][25] ),
    .B(_05171_),
    .Y(_05177_));
 sky130_fd_sc_hd__a211o_4 _10332_ (.A1(_04686_),
    .A2(_05170_),
    .B1(_05176_),
    .C1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__inv_2 _10333_ (.A(_05178_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_4 _10334_ (.A(\CPU_Dmem_value_a5[5][24] ),
    .B(_05171_),
    .Y(_05179_));
 sky130_fd_sc_hd__a211o_4 _10335_ (.A1(_04690_),
    .A2(_05170_),
    .B1(_05176_),
    .C1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__inv_2 _10336_ (.A(_05180_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_4 _10337_ (.A(\CPU_Dmem_value_a5[5][23] ),
    .B(_05171_),
    .Y(_05181_));
 sky130_fd_sc_hd__a211o_4 _10338_ (.A1(_04695_),
    .A2(_05170_),
    .B1(_05176_),
    .C1(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__inv_2 _10339_ (.A(_05182_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_4 _10340_ (.A(\CPU_Dmem_value_a5[5][22] ),
    .B(_05171_),
    .Y(_05183_));
 sky130_fd_sc_hd__a211o_4 _10341_ (.A1(_04699_),
    .A2(_05170_),
    .B1(_05176_),
    .C1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__inv_2 _10342_ (.A(_05184_),
    .Y(_01380_));
 sky130_fd_sc_hd__buf_2 _10343_ (.A(_05157_),
    .X(_05185_));
 sky130_fd_sc_hd__buf_2 _10344_ (.A(_05160_),
    .X(_05186_));
 sky130_fd_sc_hd__nor2_4 _10345_ (.A(\CPU_Dmem_value_a5[5][21] ),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__a211o_4 _10346_ (.A1(_04703_),
    .A2(_05185_),
    .B1(_05176_),
    .C1(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__inv_2 _10347_ (.A(_05188_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_4 _10348_ (.A(\CPU_Dmem_value_a5[5][20] ),
    .B(_05186_),
    .Y(_05189_));
 sky130_fd_sc_hd__a211o_4 _10349_ (.A1(_04707_),
    .A2(_05185_),
    .B1(_05176_),
    .C1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__inv_2 _10350_ (.A(_05190_),
    .Y(_01378_));
 sky130_fd_sc_hd__buf_2 _10351_ (.A(_05107_),
    .X(_05191_));
 sky130_fd_sc_hd__nor2_4 _10352_ (.A(\CPU_Dmem_value_a5[5][19] ),
    .B(_05186_),
    .Y(_05192_));
 sky130_fd_sc_hd__a211o_4 _10353_ (.A1(_04713_),
    .A2(_05185_),
    .B1(_05191_),
    .C1(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__inv_2 _10354_ (.A(_05193_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_4 _10355_ (.A(\CPU_Dmem_value_a5[5][18] ),
    .B(_05186_),
    .Y(_05194_));
 sky130_fd_sc_hd__a211o_4 _10356_ (.A1(_04717_),
    .A2(_05185_),
    .B1(_05191_),
    .C1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__inv_2 _10357_ (.A(_05195_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_4 _10358_ (.A(\CPU_Dmem_value_a5[5][17] ),
    .B(_05186_),
    .Y(_05196_));
 sky130_fd_sc_hd__a211o_4 _10359_ (.A1(_04722_),
    .A2(_05185_),
    .B1(_05191_),
    .C1(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__inv_2 _10360_ (.A(_05197_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_4 _10361_ (.A(\CPU_Dmem_value_a5[5][16] ),
    .B(_05186_),
    .Y(_05198_));
 sky130_fd_sc_hd__a211o_4 _10362_ (.A1(_04726_),
    .A2(_05185_),
    .B1(_05191_),
    .C1(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__inv_2 _10363_ (.A(_05199_),
    .Y(_01374_));
 sky130_fd_sc_hd__buf_2 _10364_ (.A(_05157_),
    .X(_05200_));
 sky130_fd_sc_hd__buf_2 _10365_ (.A(_05160_),
    .X(_05201_));
 sky130_fd_sc_hd__nor2_4 _10366_ (.A(\CPU_Dmem_value_a5[5][15] ),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__a211o_4 _10367_ (.A1(_04730_),
    .A2(_05200_),
    .B1(_05191_),
    .C1(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__inv_2 _10368_ (.A(_05203_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_4 _10369_ (.A(\CPU_Dmem_value_a5[5][14] ),
    .B(_05201_),
    .Y(_05204_));
 sky130_fd_sc_hd__a211o_4 _10370_ (.A1(_04734_),
    .A2(_05200_),
    .B1(_05191_),
    .C1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__inv_2 _10371_ (.A(_05205_),
    .Y(_01372_));
 sky130_fd_sc_hd__buf_2 _10372_ (.A(_04904_),
    .X(_05206_));
 sky130_fd_sc_hd__buf_2 _10373_ (.A(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__nor2_4 _10374_ (.A(\CPU_Dmem_value_a5[5][13] ),
    .B(_05201_),
    .Y(_05208_));
 sky130_fd_sc_hd__a211o_4 _10375_ (.A1(_04740_),
    .A2(_05200_),
    .B1(_05207_),
    .C1(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__inv_2 _10376_ (.A(_05209_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_4 _10377_ (.A(\CPU_Dmem_value_a5[5][12] ),
    .B(_05201_),
    .Y(_05210_));
 sky130_fd_sc_hd__a211o_4 _10378_ (.A1(_04744_),
    .A2(_05200_),
    .B1(_05207_),
    .C1(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__inv_2 _10379_ (.A(_05211_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_4 _10380_ (.A(\CPU_Dmem_value_a5[5][11] ),
    .B(_05201_),
    .Y(_05212_));
 sky130_fd_sc_hd__a211o_4 _10381_ (.A1(_04749_),
    .A2(_05200_),
    .B1(_05207_),
    .C1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__inv_2 _10382_ (.A(_05213_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_4 _10383_ (.A(\CPU_Dmem_value_a5[5][10] ),
    .B(_05201_),
    .Y(_05214_));
 sky130_fd_sc_hd__a211o_4 _10384_ (.A1(_04753_),
    .A2(_05200_),
    .B1(_05207_),
    .C1(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__inv_2 _10385_ (.A(_05215_),
    .Y(_01368_));
 sky130_fd_sc_hd__buf_2 _10386_ (.A(_05160_),
    .X(_05216_));
 sky130_fd_sc_hd__buf_2 _10387_ (.A(_05160_),
    .X(_05217_));
 sky130_fd_sc_hd__nor2_4 _10388_ (.A(\CPU_Dmem_value_a5[5][9] ),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__a211o_4 _10389_ (.A1(_04757_),
    .A2(_05216_),
    .B1(_05207_),
    .C1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__inv_2 _10390_ (.A(_05219_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_4 _10391_ (.A(\CPU_Dmem_value_a5[5][8] ),
    .B(_05217_),
    .Y(_05220_));
 sky130_fd_sc_hd__a211o_4 _10392_ (.A1(_04761_),
    .A2(_05216_),
    .B1(_05207_),
    .C1(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__inv_2 _10393_ (.A(_05221_),
    .Y(_01366_));
 sky130_fd_sc_hd__buf_2 _10394_ (.A(_05206_),
    .X(_05222_));
 sky130_fd_sc_hd__nor2_4 _10395_ (.A(\CPU_Dmem_value_a5[5][7] ),
    .B(_05217_),
    .Y(_05223_));
 sky130_fd_sc_hd__a211o_4 _10396_ (.A1(_04767_),
    .A2(_05216_),
    .B1(_05222_),
    .C1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__inv_2 _10397_ (.A(_05224_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_4 _10398_ (.A(\CPU_Dmem_value_a5[5][6] ),
    .B(_05217_),
    .Y(_05225_));
 sky130_fd_sc_hd__a211o_4 _10399_ (.A1(_04771_),
    .A2(_05216_),
    .B1(_05222_),
    .C1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__inv_2 _10400_ (.A(_05226_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_4 _10401_ (.A(\CPU_Dmem_value_a5[5][5] ),
    .B(_05217_),
    .Y(_05227_));
 sky130_fd_sc_hd__a211o_4 _10402_ (.A1(_04776_),
    .A2(_05216_),
    .B1(_05222_),
    .C1(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__inv_2 _10403_ (.A(_05228_),
    .Y(_01363_));
 sky130_fd_sc_hd__nor2_4 _10404_ (.A(\CPU_Dmem_value_a5[5][4] ),
    .B(_05217_),
    .Y(_05229_));
 sky130_fd_sc_hd__a211o_4 _10405_ (.A1(_04780_),
    .A2(_05216_),
    .B1(_05222_),
    .C1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__inv_2 _10406_ (.A(_05230_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_4 _10407_ (.A(\CPU_Dmem_value_a5[5][3] ),
    .B(_05157_),
    .Y(_05231_));
 sky130_fd_sc_hd__a211o_4 _10408_ (.A1(_04784_),
    .A2(_05161_),
    .B1(_05222_),
    .C1(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__inv_2 _10409_ (.A(_05232_),
    .Y(_01361_));
 sky130_fd_sc_hd__and2_4 _10410_ (.A(\CPU_Dmem_value_a5[5][2] ),
    .B(_05155_),
    .X(_05233_));
 sky130_fd_sc_hd__a211o_4 _10411_ (.A1(_05147_),
    .A2(_05158_),
    .B1(_04889_),
    .C1(_05233_),
    .X(_01360_));
 sky130_fd_sc_hd__nor2_4 _10412_ (.A(\CPU_Dmem_value_a5[5][1] ),
    .B(_05157_),
    .Y(_05234_));
 sky130_fd_sc_hd__a211o_4 _10413_ (.A1(_04794_),
    .A2(_05161_),
    .B1(_05222_),
    .C1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__inv_2 _10414_ (.A(_05235_),
    .Y(_01359_));
 sky130_fd_sc_hd__buf_2 _10415_ (.A(_04888_),
    .X(_05236_));
 sky130_fd_sc_hd__and2_4 _10416_ (.A(\CPU_Dmem_value_a5[5][0] ),
    .B(_05155_),
    .X(_05237_));
 sky130_fd_sc_hd__a211o_4 _10417_ (.A1(_04887_),
    .A2(_05158_),
    .B1(_05236_),
    .C1(_05237_),
    .X(_01358_));
 sky130_fd_sc_hd__or4_4 _10418_ (.A(_04892_),
    .B(\CPU_dmem_addr_a4[0] ),
    .C(\CPU_dmem_addr_a4[3] ),
    .D(_05066_),
    .X(_05238_));
 sky130_fd_sc_hd__buf_2 _10419_ (.A(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__nor2_4 _10420_ (.A(_04649_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__buf_2 _10421_ (.A(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__buf_2 _10422_ (.A(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__buf_2 _10423_ (.A(_05206_),
    .X(_05243_));
 sky130_fd_sc_hd__buf_2 _10424_ (.A(_05241_),
    .X(_05244_));
 sky130_fd_sc_hd__nor2_4 _10425_ (.A(\CPU_Dmem_value_a5[6][31] ),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__a211o_4 _10426_ (.A1(_04802_),
    .A2(_05242_),
    .B1(_05243_),
    .C1(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__inv_2 _10427_ (.A(_05246_),
    .Y(_01357_));
 sky130_fd_sc_hd__buf_2 _10428_ (.A(_04646_),
    .X(_05247_));
 sky130_fd_sc_hd__nor2_4 _10429_ (.A(\CPU_Dmem_value_a5[6][30] ),
    .B(_05244_),
    .Y(_05248_));
 sky130_fd_sc_hd__a211o_4 _10430_ (.A1(_05247_),
    .A2(_05242_),
    .B1(_05243_),
    .C1(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__inv_2 _10431_ (.A(_05249_),
    .Y(_01356_));
 sky130_fd_sc_hd__buf_2 _10432_ (.A(_04667_),
    .X(_05250_));
 sky130_fd_sc_hd__buf_2 _10433_ (.A(_05240_),
    .X(_05251_));
 sky130_fd_sc_hd__buf_2 _10434_ (.A(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__buf_2 _10435_ (.A(_05241_),
    .X(_05253_));
 sky130_fd_sc_hd__nor2_4 _10436_ (.A(\CPU_Dmem_value_a5[6][29] ),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a211o_4 _10437_ (.A1(_05250_),
    .A2(_05252_),
    .B1(_05243_),
    .C1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__inv_2 _10438_ (.A(_05255_),
    .Y(_01355_));
 sky130_fd_sc_hd__buf_2 _10439_ (.A(_04671_),
    .X(_05256_));
 sky130_fd_sc_hd__nor2_4 _10440_ (.A(\CPU_Dmem_value_a5[6][28] ),
    .B(_05253_),
    .Y(_05257_));
 sky130_fd_sc_hd__a211o_4 _10441_ (.A1(_05256_),
    .A2(_05252_),
    .B1(_05243_),
    .C1(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__inv_2 _10442_ (.A(_05258_),
    .Y(_01354_));
 sky130_fd_sc_hd__buf_2 _10443_ (.A(_04675_),
    .X(_05259_));
 sky130_fd_sc_hd__nor2_4 _10444_ (.A(\CPU_Dmem_value_a5[6][27] ),
    .B(_05253_),
    .Y(_05260_));
 sky130_fd_sc_hd__a211o_4 _10445_ (.A1(_05259_),
    .A2(_05252_),
    .B1(_05243_),
    .C1(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__inv_2 _10446_ (.A(_05261_),
    .Y(_01353_));
 sky130_fd_sc_hd__buf_2 _10447_ (.A(_04679_),
    .X(_05262_));
 sky130_fd_sc_hd__nor2_4 _10448_ (.A(\CPU_Dmem_value_a5[6][26] ),
    .B(_05253_),
    .Y(_05263_));
 sky130_fd_sc_hd__a211o_4 _10449_ (.A1(_05262_),
    .A2(_05252_),
    .B1(_05243_),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__inv_2 _10450_ (.A(_05264_),
    .Y(_01352_));
 sky130_fd_sc_hd__buf_2 _10451_ (.A(_04685_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_2 _10452_ (.A(_05206_),
    .X(_05266_));
 sky130_fd_sc_hd__nor2_4 _10453_ (.A(\CPU_Dmem_value_a5[6][25] ),
    .B(_05253_),
    .Y(_05267_));
 sky130_fd_sc_hd__a211o_4 _10454_ (.A1(_05265_),
    .A2(_05252_),
    .B1(_05266_),
    .C1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__inv_2 _10455_ (.A(_05268_),
    .Y(_01351_));
 sky130_fd_sc_hd__buf_2 _10456_ (.A(_04689_),
    .X(_05269_));
 sky130_fd_sc_hd__nor2_4 _10457_ (.A(\CPU_Dmem_value_a5[6][24] ),
    .B(_05253_),
    .Y(_05270_));
 sky130_fd_sc_hd__a211o_4 _10458_ (.A1(_05269_),
    .A2(_05252_),
    .B1(_05266_),
    .C1(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__inv_2 _10459_ (.A(_05271_),
    .Y(_01350_));
 sky130_fd_sc_hd__buf_2 _10460_ (.A(_04694_),
    .X(_05272_));
 sky130_fd_sc_hd__buf_2 _10461_ (.A(_05251_),
    .X(_05273_));
 sky130_fd_sc_hd__buf_2 _10462_ (.A(_05241_),
    .X(_05274_));
 sky130_fd_sc_hd__nor2_4 _10463_ (.A(\CPU_Dmem_value_a5[6][23] ),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a211o_4 _10464_ (.A1(_05272_),
    .A2(_05273_),
    .B1(_05266_),
    .C1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__inv_2 _10465_ (.A(_05276_),
    .Y(_01349_));
 sky130_fd_sc_hd__buf_2 _10466_ (.A(_04698_),
    .X(_05277_));
 sky130_fd_sc_hd__nor2_4 _10467_ (.A(\CPU_Dmem_value_a5[6][22] ),
    .B(_05274_),
    .Y(_05278_));
 sky130_fd_sc_hd__a211o_4 _10468_ (.A1(_05277_),
    .A2(_05273_),
    .B1(_05266_),
    .C1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__inv_2 _10469_ (.A(_05279_),
    .Y(_01348_));
 sky130_fd_sc_hd__buf_2 _10470_ (.A(_04702_),
    .X(_05280_));
 sky130_fd_sc_hd__nor2_4 _10471_ (.A(\CPU_Dmem_value_a5[6][21] ),
    .B(_05274_),
    .Y(_05281_));
 sky130_fd_sc_hd__a211o_4 _10472_ (.A1(_05280_),
    .A2(_05273_),
    .B1(_05266_),
    .C1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__inv_2 _10473_ (.A(_05282_),
    .Y(_01347_));
 sky130_fd_sc_hd__buf_2 _10474_ (.A(_04706_),
    .X(_05283_));
 sky130_fd_sc_hd__nor2_4 _10475_ (.A(\CPU_Dmem_value_a5[6][20] ),
    .B(_05274_),
    .Y(_05284_));
 sky130_fd_sc_hd__a211o_4 _10476_ (.A1(_05283_),
    .A2(_05273_),
    .B1(_05266_),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__inv_2 _10477_ (.A(_05285_),
    .Y(_01346_));
 sky130_fd_sc_hd__buf_2 _10478_ (.A(_04712_),
    .X(_05286_));
 sky130_fd_sc_hd__buf_2 _10479_ (.A(_05206_),
    .X(_05287_));
 sky130_fd_sc_hd__nor2_4 _10480_ (.A(\CPU_Dmem_value_a5[6][19] ),
    .B(_05274_),
    .Y(_05288_));
 sky130_fd_sc_hd__a211o_4 _10481_ (.A1(_05286_),
    .A2(_05273_),
    .B1(_05287_),
    .C1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__inv_2 _10482_ (.A(_05289_),
    .Y(_01345_));
 sky130_fd_sc_hd__buf_2 _10483_ (.A(_04716_),
    .X(_05290_));
 sky130_fd_sc_hd__nor2_4 _10484_ (.A(\CPU_Dmem_value_a5[6][18] ),
    .B(_05274_),
    .Y(_05291_));
 sky130_fd_sc_hd__a211o_4 _10485_ (.A1(_05290_),
    .A2(_05273_),
    .B1(_05287_),
    .C1(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__inv_2 _10486_ (.A(_05292_),
    .Y(_01344_));
 sky130_fd_sc_hd__buf_2 _10487_ (.A(_04721_),
    .X(_05293_));
 sky130_fd_sc_hd__buf_2 _10488_ (.A(_05241_),
    .X(_05294_));
 sky130_fd_sc_hd__buf_2 _10489_ (.A(_05240_),
    .X(_05295_));
 sky130_fd_sc_hd__nor2_4 _10490_ (.A(\CPU_Dmem_value_a5[6][17] ),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__a211o_4 _10491_ (.A1(_05293_),
    .A2(_05294_),
    .B1(_05287_),
    .C1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__inv_2 _10492_ (.A(_05297_),
    .Y(_01343_));
 sky130_fd_sc_hd__buf_2 _10493_ (.A(_04725_),
    .X(_05298_));
 sky130_fd_sc_hd__nor2_4 _10494_ (.A(\CPU_Dmem_value_a5[6][16] ),
    .B(_05295_),
    .Y(_05299_));
 sky130_fd_sc_hd__a211o_4 _10495_ (.A1(_05298_),
    .A2(_05294_),
    .B1(_05287_),
    .C1(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__inv_2 _10496_ (.A(_05300_),
    .Y(_01342_));
 sky130_fd_sc_hd__buf_2 _10497_ (.A(_04729_),
    .X(_05301_));
 sky130_fd_sc_hd__nor2_4 _10498_ (.A(\CPU_Dmem_value_a5[6][15] ),
    .B(_05295_),
    .Y(_05302_));
 sky130_fd_sc_hd__a211o_4 _10499_ (.A1(_05301_),
    .A2(_05294_),
    .B1(_05287_),
    .C1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__inv_2 _10500_ (.A(_05303_),
    .Y(_01341_));
 sky130_fd_sc_hd__buf_2 _10501_ (.A(_04733_),
    .X(_05304_));
 sky130_fd_sc_hd__nor2_4 _10502_ (.A(\CPU_Dmem_value_a5[6][14] ),
    .B(_05295_),
    .Y(_05305_));
 sky130_fd_sc_hd__a211o_4 _10503_ (.A1(_05304_),
    .A2(_05294_),
    .B1(_05287_),
    .C1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__inv_2 _10504_ (.A(_05306_),
    .Y(_01340_));
 sky130_fd_sc_hd__buf_2 _10505_ (.A(_04739_),
    .X(_05307_));
 sky130_fd_sc_hd__buf_2 _10506_ (.A(_05206_),
    .X(_05308_));
 sky130_fd_sc_hd__nor2_4 _10507_ (.A(\CPU_Dmem_value_a5[6][13] ),
    .B(_05295_),
    .Y(_05309_));
 sky130_fd_sc_hd__a211o_4 _10508_ (.A1(_05307_),
    .A2(_05294_),
    .B1(_05308_),
    .C1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__inv_2 _10509_ (.A(_05310_),
    .Y(_01339_));
 sky130_fd_sc_hd__buf_2 _10510_ (.A(_04743_),
    .X(_05311_));
 sky130_fd_sc_hd__nor2_4 _10511_ (.A(\CPU_Dmem_value_a5[6][12] ),
    .B(_05295_),
    .Y(_05312_));
 sky130_fd_sc_hd__a211o_4 _10512_ (.A1(_05311_),
    .A2(_05294_),
    .B1(_05308_),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__inv_2 _10513_ (.A(_05313_),
    .Y(_01338_));
 sky130_fd_sc_hd__buf_2 _10514_ (.A(_04748_),
    .X(_05314_));
 sky130_fd_sc_hd__buf_2 _10515_ (.A(_05241_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_2 _10516_ (.A(_05240_),
    .X(_05316_));
 sky130_fd_sc_hd__nor2_4 _10517_ (.A(\CPU_Dmem_value_a5[6][11] ),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__a211o_4 _10518_ (.A1(_05314_),
    .A2(_05315_),
    .B1(_05308_),
    .C1(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__inv_2 _10519_ (.A(_05318_),
    .Y(_01337_));
 sky130_fd_sc_hd__buf_2 _10520_ (.A(_04752_),
    .X(_05319_));
 sky130_fd_sc_hd__nor2_4 _10521_ (.A(\CPU_Dmem_value_a5[6][10] ),
    .B(_05316_),
    .Y(_05320_));
 sky130_fd_sc_hd__a211o_4 _10522_ (.A1(_05319_),
    .A2(_05315_),
    .B1(_05308_),
    .C1(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__inv_2 _10523_ (.A(_05321_),
    .Y(_01336_));
 sky130_fd_sc_hd__buf_2 _10524_ (.A(_04756_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_4 _10525_ (.A(\CPU_Dmem_value_a5[6][9] ),
    .B(_05316_),
    .Y(_05323_));
 sky130_fd_sc_hd__a211o_4 _10526_ (.A1(_05322_),
    .A2(_05315_),
    .B1(_05308_),
    .C1(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__inv_2 _10527_ (.A(_05324_),
    .Y(_01335_));
 sky130_fd_sc_hd__buf_2 _10528_ (.A(_04760_),
    .X(_05325_));
 sky130_fd_sc_hd__nor2_4 _10529_ (.A(\CPU_Dmem_value_a5[6][8] ),
    .B(_05316_),
    .Y(_05326_));
 sky130_fd_sc_hd__a211o_4 _10530_ (.A1(_05325_),
    .A2(_05315_),
    .B1(_05308_),
    .C1(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__inv_2 _10531_ (.A(_05327_),
    .Y(_01334_));
 sky130_fd_sc_hd__buf_2 _10532_ (.A(_04766_),
    .X(_05328_));
 sky130_fd_sc_hd__buf_2 _10533_ (.A(_04904_),
    .X(_05329_));
 sky130_fd_sc_hd__buf_2 _10534_ (.A(_05329_),
    .X(_05330_));
 sky130_fd_sc_hd__nor2_4 _10535_ (.A(\CPU_Dmem_value_a5[6][7] ),
    .B(_05316_),
    .Y(_05331_));
 sky130_fd_sc_hd__a211o_4 _10536_ (.A1(_05328_),
    .A2(_05315_),
    .B1(_05330_),
    .C1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__inv_2 _10537_ (.A(_05332_),
    .Y(_01333_));
 sky130_fd_sc_hd__buf_2 _10538_ (.A(_04770_),
    .X(_05333_));
 sky130_fd_sc_hd__nor2_4 _10539_ (.A(\CPU_Dmem_value_a5[6][6] ),
    .B(_05316_),
    .Y(_05334_));
 sky130_fd_sc_hd__a211o_4 _10540_ (.A1(_05333_),
    .A2(_05315_),
    .B1(_05330_),
    .C1(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__inv_2 _10541_ (.A(_05335_),
    .Y(_01332_));
 sky130_fd_sc_hd__buf_2 _10542_ (.A(_04775_),
    .X(_05336_));
 sky130_fd_sc_hd__nor2_4 _10543_ (.A(\CPU_Dmem_value_a5[6][5] ),
    .B(_05251_),
    .Y(_05337_));
 sky130_fd_sc_hd__a211o_4 _10544_ (.A1(_05336_),
    .A2(_05244_),
    .B1(_05330_),
    .C1(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__inv_2 _10545_ (.A(_05338_),
    .Y(_01331_));
 sky130_fd_sc_hd__buf_2 _10546_ (.A(_04779_),
    .X(_05339_));
 sky130_fd_sc_hd__nor2_4 _10547_ (.A(\CPU_Dmem_value_a5[6][4] ),
    .B(_05251_),
    .Y(_05340_));
 sky130_fd_sc_hd__a211o_4 _10548_ (.A1(_05339_),
    .A2(_05244_),
    .B1(_05330_),
    .C1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__inv_2 _10549_ (.A(_05341_),
    .Y(_01330_));
 sky130_fd_sc_hd__nor2_4 _10550_ (.A(\CPU_Dmem_value_a5[6][3] ),
    .B(_05251_),
    .Y(_05342_));
 sky130_fd_sc_hd__a211o_4 _10551_ (.A1(_04783_),
    .A2(_05244_),
    .B1(_05330_),
    .C1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__inv_2 _10552_ (.A(_05343_),
    .Y(_01329_));
 sky130_fd_sc_hd__inv_2 _10553_ (.A(\CPU_Dmem_value_a5[6][2] ),
    .Y(_05344_));
 sky130_fd_sc_hd__nor2_4 _10554_ (.A(_05344_),
    .B(_05242_),
    .Y(_05345_));
 sky130_fd_sc_hd__a211o_4 _10555_ (.A1(_05147_),
    .A2(_05242_),
    .B1(_05236_),
    .C1(_05345_),
    .X(_01328_));
 sky130_fd_sc_hd__inv_2 _10556_ (.A(\CPU_Dmem_value_a5[6][1] ),
    .Y(_05346_));
 sky130_fd_sc_hd__nor2_4 _10557_ (.A(_05346_),
    .B(_05242_),
    .Y(_05347_));
 sky130_fd_sc_hd__a211o_4 _10558_ (.A1(_04976_),
    .A2(_05242_),
    .B1(_05236_),
    .C1(_05347_),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_4 _10559_ (.A(\CPU_Dmem_value_a5[6][0] ),
    .B(_05251_),
    .Y(_05348_));
 sky130_fd_sc_hd__a211o_4 _10560_ (.A1(_04798_),
    .A2(_05244_),
    .B1(_05330_),
    .C1(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__inv_2 _10561_ (.A(_05349_),
    .Y(_01326_));
 sky130_fd_sc_hd__buf_2 _10562_ (.A(_04801_),
    .X(_05350_));
 sky130_fd_sc_hd__buf_2 _10563_ (.A(_04648_),
    .X(_05351_));
 sky130_fd_sc_hd__or4_4 _10564_ (.A(_04893_),
    .B(_04804_),
    .C(_04652_),
    .D(_05067_),
    .X(_05352_));
 sky130_fd_sc_hd__or2_4 _10565_ (.A(_05351_),
    .B(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__inv_2 _10566_ (.A(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__buf_2 _10567_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__buf_2 _10568_ (.A(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__buf_2 _10569_ (.A(_05329_),
    .X(_05357_));
 sky130_fd_sc_hd__buf_2 _10570_ (.A(_05354_),
    .X(_05358_));
 sky130_fd_sc_hd__nor2_4 _10571_ (.A(\CPU_Dmem_value_a5[7][31] ),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__a211o_4 _10572_ (.A1(_05350_),
    .A2(_05356_),
    .B1(_05357_),
    .C1(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__inv_2 _10573_ (.A(_05360_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_4 _10574_ (.A(\CPU_Dmem_value_a5[7][30] ),
    .B(_05358_),
    .Y(_05361_));
 sky130_fd_sc_hd__a211o_4 _10575_ (.A1(_05247_),
    .A2(_05356_),
    .B1(_05357_),
    .C1(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__inv_2 _10576_ (.A(_05362_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_4 _10577_ (.A(\CPU_Dmem_value_a5[7][29] ),
    .B(_05358_),
    .Y(_05363_));
 sky130_fd_sc_hd__a211o_4 _10578_ (.A1(_05250_),
    .A2(_05356_),
    .B1(_05357_),
    .C1(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__inv_2 _10579_ (.A(_05364_),
    .Y(_01323_));
 sky130_fd_sc_hd__buf_2 _10580_ (.A(_05355_),
    .X(_05365_));
 sky130_fd_sc_hd__nor2_4 _10581_ (.A(\CPU_Dmem_value_a5[7][28] ),
    .B(_05358_),
    .Y(_05366_));
 sky130_fd_sc_hd__a211o_4 _10582_ (.A1(_05256_),
    .A2(_05365_),
    .B1(_05357_),
    .C1(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__inv_2 _10583_ (.A(_05367_),
    .Y(_01322_));
 sky130_fd_sc_hd__buf_2 _10584_ (.A(_05354_),
    .X(_05368_));
 sky130_fd_sc_hd__nor2_4 _10585_ (.A(\CPU_Dmem_value_a5[7][27] ),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__a211o_4 _10586_ (.A1(_05259_),
    .A2(_05365_),
    .B1(_05357_),
    .C1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__inv_2 _10587_ (.A(_05370_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_4 _10588_ (.A(\CPU_Dmem_value_a5[7][26] ),
    .B(_05368_),
    .Y(_05371_));
 sky130_fd_sc_hd__a211o_4 _10589_ (.A1(_05262_),
    .A2(_05365_),
    .B1(_05357_),
    .C1(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__inv_2 _10590_ (.A(_05372_),
    .Y(_01320_));
 sky130_fd_sc_hd__buf_2 _10591_ (.A(_05329_),
    .X(_05373_));
 sky130_fd_sc_hd__nor2_4 _10592_ (.A(\CPU_Dmem_value_a5[7][25] ),
    .B(_05368_),
    .Y(_05374_));
 sky130_fd_sc_hd__a211o_4 _10593_ (.A1(_05265_),
    .A2(_05365_),
    .B1(_05373_),
    .C1(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__inv_2 _10594_ (.A(_05375_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_4 _10595_ (.A(\CPU_Dmem_value_a5[7][24] ),
    .B(_05368_),
    .Y(_05376_));
 sky130_fd_sc_hd__a211o_4 _10596_ (.A1(_05269_),
    .A2(_05365_),
    .B1(_05373_),
    .C1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__inv_2 _10597_ (.A(_05377_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_4 _10598_ (.A(\CPU_Dmem_value_a5[7][23] ),
    .B(_05368_),
    .Y(_05378_));
 sky130_fd_sc_hd__a211o_4 _10599_ (.A1(_05272_),
    .A2(_05365_),
    .B1(_05373_),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__inv_2 _10600_ (.A(_05379_),
    .Y(_01317_));
 sky130_fd_sc_hd__buf_2 _10601_ (.A(_05355_),
    .X(_05380_));
 sky130_fd_sc_hd__nor2_4 _10602_ (.A(\CPU_Dmem_value_a5[7][22] ),
    .B(_05368_),
    .Y(_05381_));
 sky130_fd_sc_hd__a211o_4 _10603_ (.A1(_05277_),
    .A2(_05380_),
    .B1(_05373_),
    .C1(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__inv_2 _10604_ (.A(_05382_),
    .Y(_01316_));
 sky130_fd_sc_hd__buf_2 _10605_ (.A(_05354_),
    .X(_05383_));
 sky130_fd_sc_hd__nor2_4 _10606_ (.A(\CPU_Dmem_value_a5[7][21] ),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__a211o_4 _10607_ (.A1(_05280_),
    .A2(_05380_),
    .B1(_05373_),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__inv_2 _10608_ (.A(_05385_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_4 _10609_ (.A(\CPU_Dmem_value_a5[7][20] ),
    .B(_05383_),
    .Y(_05386_));
 sky130_fd_sc_hd__a211o_4 _10610_ (.A1(_05283_),
    .A2(_05380_),
    .B1(_05373_),
    .C1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__inv_2 _10611_ (.A(_05387_),
    .Y(_01314_));
 sky130_fd_sc_hd__buf_2 _10612_ (.A(_05329_),
    .X(_05388_));
 sky130_fd_sc_hd__nor2_4 _10613_ (.A(\CPU_Dmem_value_a5[7][19] ),
    .B(_05383_),
    .Y(_05389_));
 sky130_fd_sc_hd__a211o_4 _10614_ (.A1(_05286_),
    .A2(_05380_),
    .B1(_05388_),
    .C1(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__inv_2 _10615_ (.A(_05390_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_4 _10616_ (.A(\CPU_Dmem_value_a5[7][18] ),
    .B(_05383_),
    .Y(_05391_));
 sky130_fd_sc_hd__a211o_4 _10617_ (.A1(_05290_),
    .A2(_05380_),
    .B1(_05388_),
    .C1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__inv_2 _10618_ (.A(_05392_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_4 _10619_ (.A(\CPU_Dmem_value_a5[7][17] ),
    .B(_05383_),
    .Y(_05393_));
 sky130_fd_sc_hd__a211o_4 _10620_ (.A1(_05293_),
    .A2(_05380_),
    .B1(_05388_),
    .C1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__inv_2 _10621_ (.A(_05394_),
    .Y(_01311_));
 sky130_fd_sc_hd__buf_2 _10622_ (.A(_05355_),
    .X(_05395_));
 sky130_fd_sc_hd__nor2_4 _10623_ (.A(\CPU_Dmem_value_a5[7][16] ),
    .B(_05383_),
    .Y(_05396_));
 sky130_fd_sc_hd__a211o_4 _10624_ (.A1(_05298_),
    .A2(_05395_),
    .B1(_05388_),
    .C1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__inv_2 _10625_ (.A(_05397_),
    .Y(_01310_));
 sky130_fd_sc_hd__buf_2 _10626_ (.A(_05354_),
    .X(_05398_));
 sky130_fd_sc_hd__nor2_4 _10627_ (.A(\CPU_Dmem_value_a5[7][15] ),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__a211o_4 _10628_ (.A1(_05301_),
    .A2(_05395_),
    .B1(_05388_),
    .C1(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__inv_2 _10629_ (.A(_05400_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_4 _10630_ (.A(\CPU_Dmem_value_a5[7][14] ),
    .B(_05398_),
    .Y(_05401_));
 sky130_fd_sc_hd__a211o_4 _10631_ (.A1(_05304_),
    .A2(_05395_),
    .B1(_05388_),
    .C1(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__inv_2 _10632_ (.A(_05402_),
    .Y(_01308_));
 sky130_fd_sc_hd__buf_2 _10633_ (.A(_05329_),
    .X(_05403_));
 sky130_fd_sc_hd__nor2_4 _10634_ (.A(\CPU_Dmem_value_a5[7][13] ),
    .B(_05398_),
    .Y(_05404_));
 sky130_fd_sc_hd__a211o_4 _10635_ (.A1(_05307_),
    .A2(_05395_),
    .B1(_05403_),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__inv_2 _10636_ (.A(_05405_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_4 _10637_ (.A(\CPU_Dmem_value_a5[7][12] ),
    .B(_05398_),
    .Y(_05406_));
 sky130_fd_sc_hd__a211o_4 _10638_ (.A1(_05311_),
    .A2(_05395_),
    .B1(_05403_),
    .C1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__inv_2 _10639_ (.A(_05407_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_4 _10640_ (.A(\CPU_Dmem_value_a5[7][11] ),
    .B(_05398_),
    .Y(_05408_));
 sky130_fd_sc_hd__a211o_4 _10641_ (.A1(_05314_),
    .A2(_05395_),
    .B1(_05403_),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__inv_2 _10642_ (.A(_05409_),
    .Y(_01305_));
 sky130_fd_sc_hd__buf_2 _10643_ (.A(_05355_),
    .X(_05410_));
 sky130_fd_sc_hd__nor2_4 _10644_ (.A(\CPU_Dmem_value_a5[7][10] ),
    .B(_05398_),
    .Y(_05411_));
 sky130_fd_sc_hd__a211o_4 _10645_ (.A1(_05319_),
    .A2(_05410_),
    .B1(_05403_),
    .C1(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__inv_2 _10646_ (.A(_05412_),
    .Y(_01304_));
 sky130_fd_sc_hd__buf_2 _10647_ (.A(_05354_),
    .X(_05413_));
 sky130_fd_sc_hd__nor2_4 _10648_ (.A(\CPU_Dmem_value_a5[7][9] ),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__a211o_4 _10649_ (.A1(_05322_),
    .A2(_05410_),
    .B1(_05403_),
    .C1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__inv_2 _10650_ (.A(_05415_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_4 _10651_ (.A(\CPU_Dmem_value_a5[7][8] ),
    .B(_05413_),
    .Y(_05416_));
 sky130_fd_sc_hd__a211o_4 _10652_ (.A1(_05325_),
    .A2(_05410_),
    .B1(_05403_),
    .C1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__inv_2 _10653_ (.A(_05417_),
    .Y(_01302_));
 sky130_fd_sc_hd__buf_2 _10654_ (.A(_05329_),
    .X(_05418_));
 sky130_fd_sc_hd__nor2_4 _10655_ (.A(\CPU_Dmem_value_a5[7][7] ),
    .B(_05413_),
    .Y(_05419_));
 sky130_fd_sc_hd__a211o_4 _10656_ (.A1(_05328_),
    .A2(_05410_),
    .B1(_05418_),
    .C1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__inv_2 _10657_ (.A(_05420_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_4 _10658_ (.A(\CPU_Dmem_value_a5[7][6] ),
    .B(_05413_),
    .Y(_05421_));
 sky130_fd_sc_hd__a211o_4 _10659_ (.A1(_05333_),
    .A2(_05410_),
    .B1(_05418_),
    .C1(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__inv_2 _10660_ (.A(_05422_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_4 _10661_ (.A(\CPU_Dmem_value_a5[7][5] ),
    .B(_05413_),
    .Y(_05423_));
 sky130_fd_sc_hd__a211o_4 _10662_ (.A1(_05336_),
    .A2(_05410_),
    .B1(_05418_),
    .C1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__inv_2 _10663_ (.A(_05424_),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2_4 _10664_ (.A(\CPU_Dmem_value_a5[7][4] ),
    .B(_05413_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211o_4 _10665_ (.A1(_05339_),
    .A2(_05358_),
    .B1(_05418_),
    .C1(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__inv_2 _10666_ (.A(_05426_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_4 _10667_ (.A(\CPU_Dmem_value_a5[7][3] ),
    .B(_05355_),
    .Y(_05427_));
 sky130_fd_sc_hd__a211o_4 _10668_ (.A1(_04783_),
    .A2(_05358_),
    .B1(_05418_),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__inv_2 _10669_ (.A(_05428_),
    .Y(_01297_));
 sky130_fd_sc_hd__and2_4 _10670_ (.A(\CPU_Dmem_value_a5[7][2] ),
    .B(_05353_),
    .X(_05429_));
 sky130_fd_sc_hd__a211o_4 _10671_ (.A1(_05147_),
    .A2(_05356_),
    .B1(_05236_),
    .C1(_05429_),
    .X(_01296_));
 sky130_fd_sc_hd__and2_4 _10672_ (.A(\CPU_Dmem_value_a5[7][1] ),
    .B(_05353_),
    .X(_05430_));
 sky130_fd_sc_hd__a211o_4 _10673_ (.A1(_04976_),
    .A2(_05356_),
    .B1(_05236_),
    .C1(_05430_),
    .X(_01295_));
 sky130_fd_sc_hd__and2_4 _10674_ (.A(\CPU_Dmem_value_a5[7][0] ),
    .B(_05353_),
    .X(_05431_));
 sky130_fd_sc_hd__a211o_4 _10675_ (.A1(_04887_),
    .A2(_05356_),
    .B1(_05236_),
    .C1(_05431_),
    .X(_01294_));
 sky130_fd_sc_hd__inv_2 _10676_ (.A(\CPU_dmem_addr_a4[3] ),
    .Y(_05432_));
 sky130_fd_sc_hd__or4_4 _10677_ (.A(\CPU_dmem_addr_a4[1] ),
    .B(\CPU_dmem_addr_a4[0] ),
    .C(_05432_),
    .D(_04653_),
    .X(_05433_));
 sky130_fd_sc_hd__buf_2 _10678_ (.A(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__nor2_4 _10679_ (.A(_04649_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__buf_2 _10680_ (.A(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__buf_2 _10681_ (.A(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__buf_2 _10682_ (.A(_05436_),
    .X(_05438_));
 sky130_fd_sc_hd__nor2_4 _10683_ (.A(\CPU_Dmem_value_a5[8][31] ),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__a211o_4 _10684_ (.A1(_05350_),
    .A2(_05437_),
    .B1(_05418_),
    .C1(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__inv_2 _10685_ (.A(_05440_),
    .Y(_01293_));
 sky130_fd_sc_hd__buf_2 _10686_ (.A(_04904_),
    .X(_05441_));
 sky130_fd_sc_hd__buf_2 _10687_ (.A(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__nor2_4 _10688_ (.A(\CPU_Dmem_value_a5[8][30] ),
    .B(_05438_),
    .Y(_05443_));
 sky130_fd_sc_hd__a211o_4 _10689_ (.A1(_05247_),
    .A2(_05437_),
    .B1(_05442_),
    .C1(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__inv_2 _10690_ (.A(_05444_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_4 _10691_ (.A(\CPU_Dmem_value_a5[8][29] ),
    .B(_05438_),
    .Y(_05445_));
 sky130_fd_sc_hd__a211o_4 _10692_ (.A1(_05250_),
    .A2(_05437_),
    .B1(_05442_),
    .C1(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__inv_2 _10693_ (.A(_05446_),
    .Y(_01291_));
 sky130_fd_sc_hd__buf_2 _10694_ (.A(_05436_),
    .X(_05447_));
 sky130_fd_sc_hd__nor2_4 _10695_ (.A(\CPU_Dmem_value_a5[8][28] ),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__a211o_4 _10696_ (.A1(_05256_),
    .A2(_05437_),
    .B1(_05442_),
    .C1(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__inv_2 _10697_ (.A(_05449_),
    .Y(_01290_));
 sky130_fd_sc_hd__buf_2 _10698_ (.A(_05435_),
    .X(_05450_));
 sky130_fd_sc_hd__buf_2 _10699_ (.A(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__nor2_4 _10700_ (.A(\CPU_Dmem_value_a5[8][27] ),
    .B(_05447_),
    .Y(_05452_));
 sky130_fd_sc_hd__a211o_4 _10701_ (.A1(_05259_),
    .A2(_05451_),
    .B1(_05442_),
    .C1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__inv_2 _10702_ (.A(_05453_),
    .Y(_01289_));
 sky130_fd_sc_hd__nor2_4 _10703_ (.A(\CPU_Dmem_value_a5[8][26] ),
    .B(_05447_),
    .Y(_05454_));
 sky130_fd_sc_hd__a211o_4 _10704_ (.A1(_05262_),
    .A2(_05451_),
    .B1(_05442_),
    .C1(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__inv_2 _10705_ (.A(_05455_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_4 _10706_ (.A(\CPU_Dmem_value_a5[8][25] ),
    .B(_05447_),
    .Y(_05456_));
 sky130_fd_sc_hd__a211o_4 _10707_ (.A1(_05265_),
    .A2(_05451_),
    .B1(_05442_),
    .C1(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__inv_2 _10708_ (.A(_05457_),
    .Y(_01287_));
 sky130_fd_sc_hd__buf_2 _10709_ (.A(_05441_),
    .X(_05458_));
 sky130_fd_sc_hd__nor2_4 _10710_ (.A(\CPU_Dmem_value_a5[8][24] ),
    .B(_05447_),
    .Y(_05459_));
 sky130_fd_sc_hd__a211o_4 _10711_ (.A1(_05269_),
    .A2(_05451_),
    .B1(_05458_),
    .C1(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__inv_2 _10712_ (.A(_05460_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_4 _10713_ (.A(\CPU_Dmem_value_a5[8][23] ),
    .B(_05447_),
    .Y(_05461_));
 sky130_fd_sc_hd__a211o_4 _10714_ (.A1(_05272_),
    .A2(_05451_),
    .B1(_05458_),
    .C1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__inv_2 _10715_ (.A(_05462_),
    .Y(_01285_));
 sky130_fd_sc_hd__buf_2 _10716_ (.A(_05436_),
    .X(_05463_));
 sky130_fd_sc_hd__nor2_4 _10717_ (.A(\CPU_Dmem_value_a5[8][22] ),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__a211o_4 _10718_ (.A1(_05277_),
    .A2(_05451_),
    .B1(_05458_),
    .C1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__inv_2 _10719_ (.A(_05465_),
    .Y(_01284_));
 sky130_fd_sc_hd__buf_2 _10720_ (.A(_05450_),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_4 _10721_ (.A(\CPU_Dmem_value_a5[8][21] ),
    .B(_05463_),
    .Y(_05467_));
 sky130_fd_sc_hd__a211o_4 _10722_ (.A1(_05280_),
    .A2(_05466_),
    .B1(_05458_),
    .C1(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__inv_2 _10723_ (.A(_05468_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_4 _10724_ (.A(\CPU_Dmem_value_a5[8][20] ),
    .B(_05463_),
    .Y(_05469_));
 sky130_fd_sc_hd__a211o_4 _10725_ (.A1(_05283_),
    .A2(_05466_),
    .B1(_05458_),
    .C1(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__inv_2 _10726_ (.A(_05470_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_4 _10727_ (.A(\CPU_Dmem_value_a5[8][19] ),
    .B(_05463_),
    .Y(_05471_));
 sky130_fd_sc_hd__a211o_4 _10728_ (.A1(_05286_),
    .A2(_05466_),
    .B1(_05458_),
    .C1(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__inv_2 _10729_ (.A(_05472_),
    .Y(_01281_));
 sky130_fd_sc_hd__buf_2 _10730_ (.A(_05441_),
    .X(_05473_));
 sky130_fd_sc_hd__nor2_4 _10731_ (.A(\CPU_Dmem_value_a5[8][18] ),
    .B(_05463_),
    .Y(_05474_));
 sky130_fd_sc_hd__a211o_4 _10732_ (.A1(_05290_),
    .A2(_05466_),
    .B1(_05473_),
    .C1(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__inv_2 _10733_ (.A(_05475_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_4 _10734_ (.A(\CPU_Dmem_value_a5[8][17] ),
    .B(_05463_),
    .Y(_05476_));
 sky130_fd_sc_hd__a211o_4 _10735_ (.A1(_05293_),
    .A2(_05466_),
    .B1(_05473_),
    .C1(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__inv_2 _10736_ (.A(_05477_),
    .Y(_01279_));
 sky130_fd_sc_hd__buf_2 _10737_ (.A(_05435_),
    .X(_05478_));
 sky130_fd_sc_hd__nor2_4 _10738_ (.A(\CPU_Dmem_value_a5[8][16] ),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__a211o_4 _10739_ (.A1(_05298_),
    .A2(_05466_),
    .B1(_05473_),
    .C1(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__inv_2 _10740_ (.A(_05480_),
    .Y(_01278_));
 sky130_fd_sc_hd__buf_2 _10741_ (.A(_05436_),
    .X(_05481_));
 sky130_fd_sc_hd__nor2_4 _10742_ (.A(\CPU_Dmem_value_a5[8][15] ),
    .B(_05478_),
    .Y(_05482_));
 sky130_fd_sc_hd__a211o_4 _10743_ (.A1(_05301_),
    .A2(_05481_),
    .B1(_05473_),
    .C1(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__inv_2 _10744_ (.A(_05483_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_4 _10745_ (.A(\CPU_Dmem_value_a5[8][14] ),
    .B(_05478_),
    .Y(_05484_));
 sky130_fd_sc_hd__a211o_4 _10746_ (.A1(_05304_),
    .A2(_05481_),
    .B1(_05473_),
    .C1(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__inv_2 _10747_ (.A(_05485_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_4 _10748_ (.A(\CPU_Dmem_value_a5[8][13] ),
    .B(_05478_),
    .Y(_05486_));
 sky130_fd_sc_hd__a211o_4 _10749_ (.A1(_05307_),
    .A2(_05481_),
    .B1(_05473_),
    .C1(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__inv_2 _10750_ (.A(_05487_),
    .Y(_01275_));
 sky130_fd_sc_hd__buf_2 _10751_ (.A(_05441_),
    .X(_05488_));
 sky130_fd_sc_hd__nor2_4 _10752_ (.A(\CPU_Dmem_value_a5[8][12] ),
    .B(_05478_),
    .Y(_05489_));
 sky130_fd_sc_hd__a211o_4 _10753_ (.A1(_05311_),
    .A2(_05481_),
    .B1(_05488_),
    .C1(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__inv_2 _10754_ (.A(_05490_),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_4 _10755_ (.A(\CPU_Dmem_value_a5[8][11] ),
    .B(_05478_),
    .Y(_05491_));
 sky130_fd_sc_hd__a211o_4 _10756_ (.A1(_05314_),
    .A2(_05481_),
    .B1(_05488_),
    .C1(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__inv_2 _10757_ (.A(_05492_),
    .Y(_01273_));
 sky130_fd_sc_hd__buf_2 _10758_ (.A(_05435_),
    .X(_05493_));
 sky130_fd_sc_hd__nor2_4 _10759_ (.A(\CPU_Dmem_value_a5[8][10] ),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__a211o_4 _10760_ (.A1(_05319_),
    .A2(_05481_),
    .B1(_05488_),
    .C1(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__inv_2 _10761_ (.A(_05495_),
    .Y(_01272_));
 sky130_fd_sc_hd__buf_2 _10762_ (.A(_05436_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_4 _10763_ (.A(\CPU_Dmem_value_a5[8][9] ),
    .B(_05493_),
    .Y(_05497_));
 sky130_fd_sc_hd__a211o_4 _10764_ (.A1(_05322_),
    .A2(_05496_),
    .B1(_05488_),
    .C1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__inv_2 _10765_ (.A(_05498_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_4 _10766_ (.A(\CPU_Dmem_value_a5[8][8] ),
    .B(_05493_),
    .Y(_05499_));
 sky130_fd_sc_hd__a211o_4 _10767_ (.A1(_05325_),
    .A2(_05496_),
    .B1(_05488_),
    .C1(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__inv_2 _10768_ (.A(_05500_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_4 _10769_ (.A(\CPU_Dmem_value_a5[8][7] ),
    .B(_05493_),
    .Y(_05501_));
 sky130_fd_sc_hd__a211o_4 _10770_ (.A1(_05328_),
    .A2(_05496_),
    .B1(_05488_),
    .C1(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__inv_2 _10771_ (.A(_05502_),
    .Y(_01269_));
 sky130_fd_sc_hd__buf_2 _10772_ (.A(_05441_),
    .X(_05503_));
 sky130_fd_sc_hd__nor2_4 _10773_ (.A(\CPU_Dmem_value_a5[8][6] ),
    .B(_05493_),
    .Y(_05504_));
 sky130_fd_sc_hd__a211o_4 _10774_ (.A1(_05333_),
    .A2(_05496_),
    .B1(_05503_),
    .C1(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__inv_2 _10775_ (.A(_05505_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_4 _10776_ (.A(\CPU_Dmem_value_a5[8][5] ),
    .B(_05493_),
    .Y(_05506_));
 sky130_fd_sc_hd__a211o_4 _10777_ (.A1(_05336_),
    .A2(_05496_),
    .B1(_05503_),
    .C1(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__inv_2 _10778_ (.A(_05507_),
    .Y(_01267_));
 sky130_fd_sc_hd__nor2_4 _10779_ (.A(\CPU_Dmem_value_a5[8][4] ),
    .B(_05450_),
    .Y(_05508_));
 sky130_fd_sc_hd__a211o_4 _10780_ (.A1(_05339_),
    .A2(_05496_),
    .B1(_05503_),
    .C1(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__inv_2 _10781_ (.A(_05509_),
    .Y(_01266_));
 sky130_fd_sc_hd__buf_2 _10782_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .X(_05510_));
 sky130_fd_sc_hd__buf_2 _10783_ (.A(_04888_),
    .X(_05511_));
 sky130_fd_sc_hd__inv_2 _10784_ (.A(\CPU_Dmem_value_a5[8][3] ),
    .Y(_05512_));
 sky130_fd_sc_hd__nor2_4 _10785_ (.A(_05512_),
    .B(_05437_),
    .Y(_05513_));
 sky130_fd_sc_hd__a211o_4 _10786_ (.A1(_05510_),
    .A2(_05437_),
    .B1(_05511_),
    .C1(_05513_),
    .X(_01265_));
 sky130_fd_sc_hd__nor2_4 _10787_ (.A(\CPU_Dmem_value_a5[8][2] ),
    .B(_05450_),
    .Y(_05514_));
 sky130_fd_sc_hd__a211o_4 _10788_ (.A1(_04788_),
    .A2(_05438_),
    .B1(_05503_),
    .C1(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__inv_2 _10789_ (.A(_05515_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_4 _10790_ (.A(\CPU_Dmem_value_a5[8][1] ),
    .B(_05450_),
    .Y(_05516_));
 sky130_fd_sc_hd__a211o_4 _10791_ (.A1(_04794_),
    .A2(_05438_),
    .B1(_05503_),
    .C1(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__inv_2 _10792_ (.A(_05517_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_4 _10793_ (.A(\CPU_Dmem_value_a5[8][0] ),
    .B(_05450_),
    .Y(_05518_));
 sky130_fd_sc_hd__a211o_4 _10794_ (.A1(_04798_),
    .A2(_05438_),
    .B1(_05503_),
    .C1(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__inv_2 _10795_ (.A(_05519_),
    .Y(_01262_));
 sky130_fd_sc_hd__or4_4 _10796_ (.A(\CPU_dmem_addr_a4[1] ),
    .B(_04803_),
    .C(_05432_),
    .D(\CPU_dmem_addr_a4[2] ),
    .X(_05520_));
 sky130_fd_sc_hd__buf_2 _10797_ (.A(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__nor2_4 _10798_ (.A(_05351_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__buf_2 _10799_ (.A(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__buf_2 _10800_ (.A(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__buf_2 _10801_ (.A(_05441_),
    .X(_05525_));
 sky130_fd_sc_hd__buf_2 _10802_ (.A(_05523_),
    .X(_05526_));
 sky130_fd_sc_hd__nor2_4 _10803_ (.A(\CPU_Dmem_value_a5[9][31] ),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a211o_4 _10804_ (.A1(_05350_),
    .A2(_05524_),
    .B1(_05525_),
    .C1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__inv_2 _10805_ (.A(_05528_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_4 _10806_ (.A(\CPU_Dmem_value_a5[9][30] ),
    .B(_05526_),
    .Y(_05529_));
 sky130_fd_sc_hd__a211o_4 _10807_ (.A1(_05247_),
    .A2(_05524_),
    .B1(_05525_),
    .C1(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__inv_2 _10808_ (.A(_05530_),
    .Y(_01260_));
 sky130_fd_sc_hd__buf_2 _10809_ (.A(_05522_),
    .X(_05531_));
 sky130_fd_sc_hd__buf_2 _10810_ (.A(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__buf_2 _10811_ (.A(_05523_),
    .X(_05533_));
 sky130_fd_sc_hd__nor2_4 _10812_ (.A(\CPU_Dmem_value_a5[9][29] ),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hd__a211o_4 _10813_ (.A1(_05250_),
    .A2(_05532_),
    .B1(_05525_),
    .C1(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__inv_2 _10814_ (.A(_05535_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_4 _10815_ (.A(\CPU_Dmem_value_a5[9][28] ),
    .B(_05533_),
    .Y(_05536_));
 sky130_fd_sc_hd__a211o_4 _10816_ (.A1(_05256_),
    .A2(_05532_),
    .B1(_05525_),
    .C1(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__inv_2 _10817_ (.A(_05537_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_4 _10818_ (.A(\CPU_Dmem_value_a5[9][27] ),
    .B(_05533_),
    .Y(_05538_));
 sky130_fd_sc_hd__a211o_4 _10819_ (.A1(_05259_),
    .A2(_05532_),
    .B1(_05525_),
    .C1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__inv_2 _10820_ (.A(_05539_),
    .Y(_01257_));
 sky130_fd_sc_hd__nor2_4 _10821_ (.A(\CPU_Dmem_value_a5[9][26] ),
    .B(_05533_),
    .Y(_05540_));
 sky130_fd_sc_hd__a211o_4 _10822_ (.A1(_05262_),
    .A2(_05532_),
    .B1(_05525_),
    .C1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__inv_2 _10823_ (.A(_05541_),
    .Y(_01256_));
 sky130_fd_sc_hd__buf_2 _10824_ (.A(_04659_),
    .X(_05542_));
 sky130_fd_sc_hd__buf_2 _10825_ (.A(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__nor2_4 _10826_ (.A(\CPU_Dmem_value_a5[9][25] ),
    .B(_05533_),
    .Y(_05544_));
 sky130_fd_sc_hd__a211o_4 _10827_ (.A1(_05265_),
    .A2(_05532_),
    .B1(_05543_),
    .C1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__inv_2 _10828_ (.A(_05545_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_4 _10829_ (.A(\CPU_Dmem_value_a5[9][24] ),
    .B(_05533_),
    .Y(_05546_));
 sky130_fd_sc_hd__a211o_4 _10830_ (.A1(_05269_),
    .A2(_05532_),
    .B1(_05543_),
    .C1(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__inv_2 _10831_ (.A(_05547_),
    .Y(_01254_));
 sky130_fd_sc_hd__buf_2 _10832_ (.A(_05531_),
    .X(_05548_));
 sky130_fd_sc_hd__buf_2 _10833_ (.A(_05523_),
    .X(_05549_));
 sky130_fd_sc_hd__nor2_4 _10834_ (.A(\CPU_Dmem_value_a5[9][23] ),
    .B(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a211o_4 _10835_ (.A1(_05272_),
    .A2(_05548_),
    .B1(_05543_),
    .C1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__inv_2 _10836_ (.A(_05551_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_4 _10837_ (.A(\CPU_Dmem_value_a5[9][22] ),
    .B(_05549_),
    .Y(_05552_));
 sky130_fd_sc_hd__a211o_4 _10838_ (.A1(_05277_),
    .A2(_05548_),
    .B1(_05543_),
    .C1(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__inv_2 _10839_ (.A(_05553_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_4 _10840_ (.A(\CPU_Dmem_value_a5[9][21] ),
    .B(_05549_),
    .Y(_05554_));
 sky130_fd_sc_hd__a211o_4 _10841_ (.A1(_05280_),
    .A2(_05548_),
    .B1(_05543_),
    .C1(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__inv_2 _10842_ (.A(_05555_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_4 _10843_ (.A(\CPU_Dmem_value_a5[9][20] ),
    .B(_05549_),
    .Y(_05556_));
 sky130_fd_sc_hd__a211o_4 _10844_ (.A1(_05283_),
    .A2(_05548_),
    .B1(_05543_),
    .C1(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__inv_2 _10845_ (.A(_05557_),
    .Y(_01250_));
 sky130_fd_sc_hd__buf_2 _10846_ (.A(_05542_),
    .X(_05558_));
 sky130_fd_sc_hd__nor2_4 _10847_ (.A(\CPU_Dmem_value_a5[9][19] ),
    .B(_05549_),
    .Y(_05559_));
 sky130_fd_sc_hd__a211o_4 _10848_ (.A1(_05286_),
    .A2(_05548_),
    .B1(_05558_),
    .C1(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__inv_2 _10849_ (.A(_05560_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_4 _10850_ (.A(\CPU_Dmem_value_a5[9][18] ),
    .B(_05549_),
    .Y(_05561_));
 sky130_fd_sc_hd__a211o_4 _10851_ (.A1(_05290_),
    .A2(_05548_),
    .B1(_05558_),
    .C1(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__inv_2 _10852_ (.A(_05562_),
    .Y(_01248_));
 sky130_fd_sc_hd__buf_2 _10853_ (.A(_05523_),
    .X(_05563_));
 sky130_fd_sc_hd__buf_2 _10854_ (.A(_05522_),
    .X(_05564_));
 sky130_fd_sc_hd__nor2_4 _10855_ (.A(\CPU_Dmem_value_a5[9][17] ),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__a211o_4 _10856_ (.A1(_05293_),
    .A2(_05563_),
    .B1(_05558_),
    .C1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__inv_2 _10857_ (.A(_05566_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_4 _10858_ (.A(\CPU_Dmem_value_a5[9][16] ),
    .B(_05564_),
    .Y(_05567_));
 sky130_fd_sc_hd__a211o_4 _10859_ (.A1(_05298_),
    .A2(_05563_),
    .B1(_05558_),
    .C1(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__inv_2 _10860_ (.A(_05568_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_4 _10861_ (.A(\CPU_Dmem_value_a5[9][15] ),
    .B(_05564_),
    .Y(_05569_));
 sky130_fd_sc_hd__a211o_4 _10862_ (.A1(_05301_),
    .A2(_05563_),
    .B1(_05558_),
    .C1(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__inv_2 _10863_ (.A(_05570_),
    .Y(_01245_));
 sky130_fd_sc_hd__nor2_4 _10864_ (.A(\CPU_Dmem_value_a5[9][14] ),
    .B(_05564_),
    .Y(_05571_));
 sky130_fd_sc_hd__a211o_4 _10865_ (.A1(_05304_),
    .A2(_05563_),
    .B1(_05558_),
    .C1(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__inv_2 _10866_ (.A(_05572_),
    .Y(_01244_));
 sky130_fd_sc_hd__buf_2 _10867_ (.A(_05542_),
    .X(_05573_));
 sky130_fd_sc_hd__nor2_4 _10868_ (.A(\CPU_Dmem_value_a5[9][13] ),
    .B(_05564_),
    .Y(_05574_));
 sky130_fd_sc_hd__a211o_4 _10869_ (.A1(_05307_),
    .A2(_05563_),
    .B1(_05573_),
    .C1(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__inv_2 _10870_ (.A(_05575_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_4 _10871_ (.A(\CPU_Dmem_value_a5[9][12] ),
    .B(_05564_),
    .Y(_05576_));
 sky130_fd_sc_hd__a211o_4 _10872_ (.A1(_05311_),
    .A2(_05563_),
    .B1(_05573_),
    .C1(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__inv_2 _10873_ (.A(_05577_),
    .Y(_01242_));
 sky130_fd_sc_hd__buf_2 _10874_ (.A(_05523_),
    .X(_05578_));
 sky130_fd_sc_hd__buf_2 _10875_ (.A(_05522_),
    .X(_05579_));
 sky130_fd_sc_hd__nor2_4 _10876_ (.A(\CPU_Dmem_value_a5[9][11] ),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a211o_4 _10877_ (.A1(_05314_),
    .A2(_05578_),
    .B1(_05573_),
    .C1(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__inv_2 _10878_ (.A(_05581_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_4 _10879_ (.A(\CPU_Dmem_value_a5[9][10] ),
    .B(_05579_),
    .Y(_05582_));
 sky130_fd_sc_hd__a211o_4 _10880_ (.A1(_05319_),
    .A2(_05578_),
    .B1(_05573_),
    .C1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__inv_2 _10881_ (.A(_05583_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_4 _10882_ (.A(\CPU_Dmem_value_a5[9][9] ),
    .B(_05579_),
    .Y(_05584_));
 sky130_fd_sc_hd__a211o_4 _10883_ (.A1(_05322_),
    .A2(_05578_),
    .B1(_05573_),
    .C1(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__inv_2 _10884_ (.A(_05585_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_4 _10885_ (.A(\CPU_Dmem_value_a5[9][8] ),
    .B(_05579_),
    .Y(_05586_));
 sky130_fd_sc_hd__a211o_4 _10886_ (.A1(_05325_),
    .A2(_05578_),
    .B1(_05573_),
    .C1(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__inv_2 _10887_ (.A(_05587_),
    .Y(_01238_));
 sky130_fd_sc_hd__buf_2 _10888_ (.A(_05542_),
    .X(_05588_));
 sky130_fd_sc_hd__nor2_4 _10889_ (.A(\CPU_Dmem_value_a5[9][7] ),
    .B(_05579_),
    .Y(_05589_));
 sky130_fd_sc_hd__a211o_4 _10890_ (.A1(_05328_),
    .A2(_05578_),
    .B1(_05588_),
    .C1(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__inv_2 _10891_ (.A(_05590_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_4 _10892_ (.A(\CPU_Dmem_value_a5[9][6] ),
    .B(_05579_),
    .Y(_05591_));
 sky130_fd_sc_hd__a211o_4 _10893_ (.A1(_05333_),
    .A2(_05578_),
    .B1(_05588_),
    .C1(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__inv_2 _10894_ (.A(_05592_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_4 _10895_ (.A(\CPU_Dmem_value_a5[9][5] ),
    .B(_05531_),
    .Y(_05593_));
 sky130_fd_sc_hd__a211o_4 _10896_ (.A1(_05336_),
    .A2(_05526_),
    .B1(_05588_),
    .C1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__inv_2 _10897_ (.A(_05594_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor2_4 _10898_ (.A(\CPU_Dmem_value_a5[9][4] ),
    .B(_05531_),
    .Y(_05595_));
 sky130_fd_sc_hd__a211o_4 _10899_ (.A1(_05339_),
    .A2(_05526_),
    .B1(_05588_),
    .C1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__inv_2 _10900_ (.A(_05596_),
    .Y(_01234_));
 sky130_fd_sc_hd__inv_2 _10901_ (.A(\CPU_Dmem_value_a5[9][3] ),
    .Y(_05597_));
 sky130_fd_sc_hd__nor2_4 _10902_ (.A(_05597_),
    .B(_05524_),
    .Y(_05598_));
 sky130_fd_sc_hd__a211o_4 _10903_ (.A1(_05510_),
    .A2(_05524_),
    .B1(_05511_),
    .C1(_05598_),
    .X(_01233_));
 sky130_fd_sc_hd__nor2_4 _10904_ (.A(\CPU_Dmem_value_a5[9][2] ),
    .B(_05531_),
    .Y(_05599_));
 sky130_fd_sc_hd__a211o_4 _10905_ (.A1(_04788_),
    .A2(_05526_),
    .B1(_05588_),
    .C1(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__inv_2 _10906_ (.A(_05600_),
    .Y(_01232_));
 sky130_fd_sc_hd__nor2_4 _10907_ (.A(\CPU_Dmem_value_a5[9][1] ),
    .B(_05531_),
    .Y(_05601_));
 sky130_fd_sc_hd__a211o_4 _10908_ (.A1(_04794_),
    .A2(_05526_),
    .B1(_05588_),
    .C1(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__inv_2 _10909_ (.A(_05602_),
    .Y(_01231_));
 sky130_fd_sc_hd__inv_2 _10910_ (.A(\CPU_Dmem_value_a5[9][0] ),
    .Y(_05603_));
 sky130_fd_sc_hd__nor2_4 _10911_ (.A(_05603_),
    .B(_05524_),
    .Y(_05604_));
 sky130_fd_sc_hd__a211o_4 _10912_ (.A1(_04887_),
    .A2(_05524_),
    .B1(_05511_),
    .C1(_05604_),
    .X(_01230_));
 sky130_fd_sc_hd__buf_2 _10913_ (.A(_05432_),
    .X(_05605_));
 sky130_fd_sc_hd__or4_4 _10914_ (.A(_04893_),
    .B(_04651_),
    .C(_05605_),
    .D(_04653_),
    .X(_05606_));
 sky130_fd_sc_hd__or2_4 _10915_ (.A(_04648_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__inv_2 _10916_ (.A(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__buf_2 _10917_ (.A(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_2 _10918_ (.A(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__buf_2 _10919_ (.A(_05542_),
    .X(_05611_));
 sky130_fd_sc_hd__buf_2 _10920_ (.A(_05608_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_2 _10921_ (.A(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__nor2_4 _10922_ (.A(\CPU_Dmem_value_a5[10][31] ),
    .B(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__a211o_4 _10923_ (.A1(_05350_),
    .A2(_05610_),
    .B1(_05611_),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__inv_2 _10924_ (.A(_05615_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_4 _10925_ (.A(\CPU_Dmem_value_a5[10][30] ),
    .B(_05613_),
    .Y(_05616_));
 sky130_fd_sc_hd__a211o_4 _10926_ (.A1(_05247_),
    .A2(_05610_),
    .B1(_05611_),
    .C1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__inv_2 _10927_ (.A(_05617_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_4 _10928_ (.A(\CPU_Dmem_value_a5[10][29] ),
    .B(_05613_),
    .Y(_05618_));
 sky130_fd_sc_hd__a211o_4 _10929_ (.A1(_05250_),
    .A2(_05610_),
    .B1(_05611_),
    .C1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__inv_2 _10930_ (.A(_05619_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_4 _10931_ (.A(\CPU_Dmem_value_a5[10][28] ),
    .B(_05613_),
    .Y(_05620_));
 sky130_fd_sc_hd__a211o_4 _10932_ (.A1(_05256_),
    .A2(_05610_),
    .B1(_05611_),
    .C1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__inv_2 _10933_ (.A(_05621_),
    .Y(_01226_));
 sky130_fd_sc_hd__buf_2 _10934_ (.A(_05609_),
    .X(_05622_));
 sky130_fd_sc_hd__buf_2 _10935_ (.A(_05612_),
    .X(_05623_));
 sky130_fd_sc_hd__nor2_4 _10936_ (.A(\CPU_Dmem_value_a5[10][27] ),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__a211o_4 _10937_ (.A1(_05259_),
    .A2(_05622_),
    .B1(_05611_),
    .C1(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__inv_2 _10938_ (.A(_05625_),
    .Y(_01225_));
 sky130_fd_sc_hd__nor2_4 _10939_ (.A(\CPU_Dmem_value_a5[10][26] ),
    .B(_05623_),
    .Y(_05626_));
 sky130_fd_sc_hd__a211o_4 _10940_ (.A1(_05262_),
    .A2(_05622_),
    .B1(_05611_),
    .C1(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__inv_2 _10941_ (.A(_05627_),
    .Y(_01224_));
 sky130_fd_sc_hd__buf_2 _10942_ (.A(_05542_),
    .X(_05628_));
 sky130_fd_sc_hd__nor2_4 _10943_ (.A(\CPU_Dmem_value_a5[10][25] ),
    .B(_05623_),
    .Y(_05629_));
 sky130_fd_sc_hd__a211o_4 _10944_ (.A1(_05265_),
    .A2(_05622_),
    .B1(_05628_),
    .C1(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__inv_2 _10945_ (.A(_05630_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_4 _10946_ (.A(\CPU_Dmem_value_a5[10][24] ),
    .B(_05623_),
    .Y(_05631_));
 sky130_fd_sc_hd__a211o_4 _10947_ (.A1(_05269_),
    .A2(_05622_),
    .B1(_05628_),
    .C1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__inv_2 _10948_ (.A(_05632_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_4 _10949_ (.A(\CPU_Dmem_value_a5[10][23] ),
    .B(_05623_),
    .Y(_05633_));
 sky130_fd_sc_hd__a211o_4 _10950_ (.A1(_05272_),
    .A2(_05622_),
    .B1(_05628_),
    .C1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__inv_2 _10951_ (.A(_05634_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_4 _10952_ (.A(\CPU_Dmem_value_a5[10][22] ),
    .B(_05623_),
    .Y(_05635_));
 sky130_fd_sc_hd__a211o_4 _10953_ (.A1(_05277_),
    .A2(_05622_),
    .B1(_05628_),
    .C1(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__inv_2 _10954_ (.A(_05636_),
    .Y(_01220_));
 sky130_fd_sc_hd__buf_2 _10955_ (.A(_05609_),
    .X(_05637_));
 sky130_fd_sc_hd__buf_2 _10956_ (.A(_05612_),
    .X(_05638_));
 sky130_fd_sc_hd__nor2_4 _10957_ (.A(\CPU_Dmem_value_a5[10][21] ),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a211o_4 _10958_ (.A1(_05280_),
    .A2(_05637_),
    .B1(_05628_),
    .C1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__inv_2 _10959_ (.A(_05640_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_4 _10960_ (.A(\CPU_Dmem_value_a5[10][20] ),
    .B(_05638_),
    .Y(_05641_));
 sky130_fd_sc_hd__a211o_4 _10961_ (.A1(_05283_),
    .A2(_05637_),
    .B1(_05628_),
    .C1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__inv_2 _10962_ (.A(_05642_),
    .Y(_01218_));
 sky130_fd_sc_hd__buf_2 _10963_ (.A(_04659_),
    .X(_05643_));
 sky130_fd_sc_hd__buf_2 _10964_ (.A(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__nor2_4 _10965_ (.A(\CPU_Dmem_value_a5[10][19] ),
    .B(_05638_),
    .Y(_05645_));
 sky130_fd_sc_hd__a211o_4 _10966_ (.A1(_05286_),
    .A2(_05637_),
    .B1(_05644_),
    .C1(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__inv_2 _10967_ (.A(_05646_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_4 _10968_ (.A(\CPU_Dmem_value_a5[10][18] ),
    .B(_05638_),
    .Y(_05647_));
 sky130_fd_sc_hd__a211o_4 _10969_ (.A1(_05290_),
    .A2(_05637_),
    .B1(_05644_),
    .C1(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__inv_2 _10970_ (.A(_05648_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_4 _10971_ (.A(\CPU_Dmem_value_a5[10][17] ),
    .B(_05638_),
    .Y(_05649_));
 sky130_fd_sc_hd__a211o_4 _10972_ (.A1(_05293_),
    .A2(_05637_),
    .B1(_05644_),
    .C1(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__inv_2 _10973_ (.A(_05650_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_4 _10974_ (.A(\CPU_Dmem_value_a5[10][16] ),
    .B(_05638_),
    .Y(_05651_));
 sky130_fd_sc_hd__a211o_4 _10975_ (.A1(_05298_),
    .A2(_05637_),
    .B1(_05644_),
    .C1(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__inv_2 _10976_ (.A(_05652_),
    .Y(_01214_));
 sky130_fd_sc_hd__buf_2 _10977_ (.A(_05609_),
    .X(_05653_));
 sky130_fd_sc_hd__buf_2 _10978_ (.A(_05612_),
    .X(_05654_));
 sky130_fd_sc_hd__nor2_4 _10979_ (.A(\CPU_Dmem_value_a5[10][15] ),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__a211o_4 _10980_ (.A1(_05301_),
    .A2(_05653_),
    .B1(_05644_),
    .C1(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__inv_2 _10981_ (.A(_05656_),
    .Y(_01213_));
 sky130_fd_sc_hd__nor2_4 _10982_ (.A(\CPU_Dmem_value_a5[10][14] ),
    .B(_05654_),
    .Y(_05657_));
 sky130_fd_sc_hd__a211o_4 _10983_ (.A1(_05304_),
    .A2(_05653_),
    .B1(_05644_),
    .C1(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__inv_2 _10984_ (.A(_05658_),
    .Y(_01212_));
 sky130_fd_sc_hd__buf_2 _10985_ (.A(_05643_),
    .X(_05659_));
 sky130_fd_sc_hd__nor2_4 _10986_ (.A(\CPU_Dmem_value_a5[10][13] ),
    .B(_05654_),
    .Y(_05660_));
 sky130_fd_sc_hd__a211o_4 _10987_ (.A1(_05307_),
    .A2(_05653_),
    .B1(_05659_),
    .C1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__inv_2 _10988_ (.A(_05661_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_4 _10989_ (.A(\CPU_Dmem_value_a5[10][12] ),
    .B(_05654_),
    .Y(_05662_));
 sky130_fd_sc_hd__a211o_4 _10990_ (.A1(_05311_),
    .A2(_05653_),
    .B1(_05659_),
    .C1(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__inv_2 _10991_ (.A(_05663_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_4 _10992_ (.A(\CPU_Dmem_value_a5[10][11] ),
    .B(_05654_),
    .Y(_05664_));
 sky130_fd_sc_hd__a211o_4 _10993_ (.A1(_05314_),
    .A2(_05653_),
    .B1(_05659_),
    .C1(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__inv_2 _10994_ (.A(_05665_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_4 _10995_ (.A(\CPU_Dmem_value_a5[10][10] ),
    .B(_05654_),
    .Y(_05666_));
 sky130_fd_sc_hd__a211o_4 _10996_ (.A1(_05319_),
    .A2(_05653_),
    .B1(_05659_),
    .C1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__inv_2 _10997_ (.A(_05667_),
    .Y(_01208_));
 sky130_fd_sc_hd__buf_2 _10998_ (.A(_05612_),
    .X(_05668_));
 sky130_fd_sc_hd__buf_2 _10999_ (.A(_05612_),
    .X(_05669_));
 sky130_fd_sc_hd__nor2_4 _11000_ (.A(\CPU_Dmem_value_a5[10][9] ),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__a211o_4 _11001_ (.A1(_05322_),
    .A2(_05668_),
    .B1(_05659_),
    .C1(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__inv_2 _11002_ (.A(_05671_),
    .Y(_01207_));
 sky130_fd_sc_hd__nor2_4 _11003_ (.A(\CPU_Dmem_value_a5[10][8] ),
    .B(_05669_),
    .Y(_05672_));
 sky130_fd_sc_hd__a211o_4 _11004_ (.A1(_05325_),
    .A2(_05668_),
    .B1(_05659_),
    .C1(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__inv_2 _11005_ (.A(_05673_),
    .Y(_01206_));
 sky130_fd_sc_hd__buf_2 _11006_ (.A(_05643_),
    .X(_05674_));
 sky130_fd_sc_hd__nor2_4 _11007_ (.A(\CPU_Dmem_value_a5[10][7] ),
    .B(_05669_),
    .Y(_05675_));
 sky130_fd_sc_hd__a211o_4 _11008_ (.A1(_05328_),
    .A2(_05668_),
    .B1(_05674_),
    .C1(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__inv_2 _11009_ (.A(_05676_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_4 _11010_ (.A(\CPU_Dmem_value_a5[10][6] ),
    .B(_05669_),
    .Y(_05677_));
 sky130_fd_sc_hd__a211o_4 _11011_ (.A1(_05333_),
    .A2(_05668_),
    .B1(_05674_),
    .C1(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__inv_2 _11012_ (.A(_05678_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_4 _11013_ (.A(\CPU_Dmem_value_a5[10][5] ),
    .B(_05669_),
    .Y(_05679_));
 sky130_fd_sc_hd__a211o_4 _11014_ (.A1(_05336_),
    .A2(_05668_),
    .B1(_05674_),
    .C1(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__inv_2 _11015_ (.A(_05680_),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_4 _11016_ (.A(\CPU_Dmem_value_a5[10][4] ),
    .B(_05669_),
    .Y(_05681_));
 sky130_fd_sc_hd__a211o_4 _11017_ (.A1(_05339_),
    .A2(_05668_),
    .B1(_05674_),
    .C1(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__inv_2 _11018_ (.A(_05682_),
    .Y(_01202_));
 sky130_fd_sc_hd__and2_4 _11019_ (.A(\CPU_Dmem_value_a5[10][3] ),
    .B(_05607_),
    .X(_05683_));
 sky130_fd_sc_hd__a211o_4 _11020_ (.A1(_05510_),
    .A2(_05610_),
    .B1(_05511_),
    .C1(_05683_),
    .X(_01201_));
 sky130_fd_sc_hd__nor2_4 _11021_ (.A(\CPU_Dmem_value_a5[10][2] ),
    .B(_05609_),
    .Y(_05684_));
 sky130_fd_sc_hd__a211o_4 _11022_ (.A1(_04787_),
    .A2(_05613_),
    .B1(_05674_),
    .C1(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__inv_2 _11023_ (.A(_05685_),
    .Y(_01200_));
 sky130_fd_sc_hd__and2_4 _11024_ (.A(\CPU_Dmem_value_a5[10][1] ),
    .B(_05607_),
    .X(_05686_));
 sky130_fd_sc_hd__a211o_4 _11025_ (.A1(_04976_),
    .A2(_05610_),
    .B1(_05511_),
    .C1(_05686_),
    .X(_01199_));
 sky130_fd_sc_hd__nor2_4 _11026_ (.A(\CPU_Dmem_value_a5[10][0] ),
    .B(_05609_),
    .Y(_05687_));
 sky130_fd_sc_hd__a211o_4 _11027_ (.A1(_04798_),
    .A2(_05613_),
    .B1(_05674_),
    .C1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__inv_2 _11028_ (.A(_05688_),
    .Y(_01198_));
 sky130_fd_sc_hd__or4_4 _11029_ (.A(_04893_),
    .B(_04804_),
    .C(_05605_),
    .D(_04653_),
    .X(_05689_));
 sky130_fd_sc_hd__or2_4 _11030_ (.A(_05351_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__inv_2 _11031_ (.A(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__buf_2 _11032_ (.A(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__buf_2 _11033_ (.A(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__buf_2 _11034_ (.A(_05643_),
    .X(_05694_));
 sky130_fd_sc_hd__buf_2 _11035_ (.A(_05691_),
    .X(_05695_));
 sky130_fd_sc_hd__nor2_4 _11036_ (.A(\CPU_Dmem_value_a5[11][31] ),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__a211o_4 _11037_ (.A1(_05350_),
    .A2(_05693_),
    .B1(_05694_),
    .C1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__inv_2 _11038_ (.A(_05697_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_4 _11039_ (.A(\CPU_Dmem_value_a5[11][30] ),
    .B(_05695_),
    .Y(_05698_));
 sky130_fd_sc_hd__a211o_4 _11040_ (.A1(_05247_),
    .A2(_05693_),
    .B1(_05694_),
    .C1(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__inv_2 _11041_ (.A(_05699_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_4 _11042_ (.A(\CPU_Dmem_value_a5[11][29] ),
    .B(_05695_),
    .Y(_05700_));
 sky130_fd_sc_hd__a211o_4 _11043_ (.A1(_05250_),
    .A2(_05693_),
    .B1(_05694_),
    .C1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__inv_2 _11044_ (.A(_05701_),
    .Y(_01195_));
 sky130_fd_sc_hd__buf_2 _11045_ (.A(_05692_),
    .X(_05702_));
 sky130_fd_sc_hd__nor2_4 _11046_ (.A(\CPU_Dmem_value_a5[11][28] ),
    .B(_05695_),
    .Y(_05703_));
 sky130_fd_sc_hd__a211o_4 _11047_ (.A1(_05256_),
    .A2(_05702_),
    .B1(_05694_),
    .C1(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__inv_2 _11048_ (.A(_05704_),
    .Y(_01194_));
 sky130_fd_sc_hd__buf_2 _11049_ (.A(_05691_),
    .X(_05705_));
 sky130_fd_sc_hd__nor2_4 _11050_ (.A(\CPU_Dmem_value_a5[11][27] ),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__a211o_4 _11051_ (.A1(_05259_),
    .A2(_05702_),
    .B1(_05694_),
    .C1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__inv_2 _11052_ (.A(_05707_),
    .Y(_01193_));
 sky130_fd_sc_hd__nor2_4 _11053_ (.A(\CPU_Dmem_value_a5[11][26] ),
    .B(_05705_),
    .Y(_05708_));
 sky130_fd_sc_hd__a211o_4 _11054_ (.A1(_05262_),
    .A2(_05702_),
    .B1(_05694_),
    .C1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__inv_2 _11055_ (.A(_05709_),
    .Y(_01192_));
 sky130_fd_sc_hd__buf_2 _11056_ (.A(_05643_),
    .X(_05710_));
 sky130_fd_sc_hd__nor2_4 _11057_ (.A(\CPU_Dmem_value_a5[11][25] ),
    .B(_05705_),
    .Y(_05711_));
 sky130_fd_sc_hd__a211o_4 _11058_ (.A1(_05265_),
    .A2(_05702_),
    .B1(_05710_),
    .C1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__inv_2 _11059_ (.A(_05712_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_4 _11060_ (.A(\CPU_Dmem_value_a5[11][24] ),
    .B(_05705_),
    .Y(_05713_));
 sky130_fd_sc_hd__a211o_4 _11061_ (.A1(_05269_),
    .A2(_05702_),
    .B1(_05710_),
    .C1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__inv_2 _11062_ (.A(_05714_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_4 _11063_ (.A(\CPU_Dmem_value_a5[11][23] ),
    .B(_05705_),
    .Y(_05715_));
 sky130_fd_sc_hd__a211o_4 _11064_ (.A1(_05272_),
    .A2(_05702_),
    .B1(_05710_),
    .C1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__inv_2 _11065_ (.A(_05716_),
    .Y(_01189_));
 sky130_fd_sc_hd__buf_2 _11066_ (.A(_05692_),
    .X(_05717_));
 sky130_fd_sc_hd__nor2_4 _11067_ (.A(\CPU_Dmem_value_a5[11][22] ),
    .B(_05705_),
    .Y(_05718_));
 sky130_fd_sc_hd__a211o_4 _11068_ (.A1(_05277_),
    .A2(_05717_),
    .B1(_05710_),
    .C1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__inv_2 _11069_ (.A(_05719_),
    .Y(_01188_));
 sky130_fd_sc_hd__buf_2 _11070_ (.A(_05691_),
    .X(_05720_));
 sky130_fd_sc_hd__nor2_4 _11071_ (.A(\CPU_Dmem_value_a5[11][21] ),
    .B(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__a211o_4 _11072_ (.A1(_05280_),
    .A2(_05717_),
    .B1(_05710_),
    .C1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__inv_2 _11073_ (.A(_05722_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_4 _11074_ (.A(\CPU_Dmem_value_a5[11][20] ),
    .B(_05720_),
    .Y(_05723_));
 sky130_fd_sc_hd__a211o_4 _11075_ (.A1(_05283_),
    .A2(_05717_),
    .B1(_05710_),
    .C1(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__inv_2 _11076_ (.A(_05724_),
    .Y(_01186_));
 sky130_fd_sc_hd__buf_2 _11077_ (.A(_05643_),
    .X(_05725_));
 sky130_fd_sc_hd__nor2_4 _11078_ (.A(\CPU_Dmem_value_a5[11][19] ),
    .B(_05720_),
    .Y(_05726_));
 sky130_fd_sc_hd__a211o_4 _11079_ (.A1(_05286_),
    .A2(_05717_),
    .B1(_05725_),
    .C1(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__inv_2 _11080_ (.A(_05727_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_4 _11081_ (.A(\CPU_Dmem_value_a5[11][18] ),
    .B(_05720_),
    .Y(_05728_));
 sky130_fd_sc_hd__a211o_4 _11082_ (.A1(_05290_),
    .A2(_05717_),
    .B1(_05725_),
    .C1(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__inv_2 _11083_ (.A(_05729_),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_4 _11084_ (.A(\CPU_Dmem_value_a5[11][17] ),
    .B(_05720_),
    .Y(_05730_));
 sky130_fd_sc_hd__a211o_4 _11085_ (.A1(_05293_),
    .A2(_05717_),
    .B1(_05725_),
    .C1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__inv_2 _11086_ (.A(_05731_),
    .Y(_01183_));
 sky130_fd_sc_hd__buf_2 _11087_ (.A(_05692_),
    .X(_05732_));
 sky130_fd_sc_hd__nor2_4 _11088_ (.A(\CPU_Dmem_value_a5[11][16] ),
    .B(_05720_),
    .Y(_05733_));
 sky130_fd_sc_hd__a211o_4 _11089_ (.A1(_05298_),
    .A2(_05732_),
    .B1(_05725_),
    .C1(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__inv_2 _11090_ (.A(_05734_),
    .Y(_01182_));
 sky130_fd_sc_hd__buf_2 _11091_ (.A(_05691_),
    .X(_05735_));
 sky130_fd_sc_hd__nor2_4 _11092_ (.A(\CPU_Dmem_value_a5[11][15] ),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__a211o_4 _11093_ (.A1(_05301_),
    .A2(_05732_),
    .B1(_05725_),
    .C1(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__inv_2 _11094_ (.A(_05737_),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2_4 _11095_ (.A(\CPU_Dmem_value_a5[11][14] ),
    .B(_05735_),
    .Y(_05738_));
 sky130_fd_sc_hd__a211o_4 _11096_ (.A1(_05304_),
    .A2(_05732_),
    .B1(_05725_),
    .C1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__inv_2 _11097_ (.A(_05739_),
    .Y(_01180_));
 sky130_fd_sc_hd__buf_2 _11098_ (.A(_04659_),
    .X(_05740_));
 sky130_fd_sc_hd__buf_2 _11099_ (.A(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__nor2_4 _11100_ (.A(\CPU_Dmem_value_a5[11][13] ),
    .B(_05735_),
    .Y(_05742_));
 sky130_fd_sc_hd__a211o_4 _11101_ (.A1(_05307_),
    .A2(_05732_),
    .B1(_05741_),
    .C1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__inv_2 _11102_ (.A(_05743_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_4 _11103_ (.A(\CPU_Dmem_value_a5[11][12] ),
    .B(_05735_),
    .Y(_05744_));
 sky130_fd_sc_hd__a211o_4 _11104_ (.A1(_05311_),
    .A2(_05732_),
    .B1(_05741_),
    .C1(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__inv_2 _11105_ (.A(_05745_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor2_4 _11106_ (.A(\CPU_Dmem_value_a5[11][11] ),
    .B(_05735_),
    .Y(_05746_));
 sky130_fd_sc_hd__a211o_4 _11107_ (.A1(_05314_),
    .A2(_05732_),
    .B1(_05741_),
    .C1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__inv_2 _11108_ (.A(_05747_),
    .Y(_01177_));
 sky130_fd_sc_hd__buf_2 _11109_ (.A(_05692_),
    .X(_05748_));
 sky130_fd_sc_hd__nor2_4 _11110_ (.A(\CPU_Dmem_value_a5[11][10] ),
    .B(_05735_),
    .Y(_05749_));
 sky130_fd_sc_hd__a211o_4 _11111_ (.A1(_05319_),
    .A2(_05748_),
    .B1(_05741_),
    .C1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__inv_2 _11112_ (.A(_05750_),
    .Y(_01176_));
 sky130_fd_sc_hd__buf_2 _11113_ (.A(_05691_),
    .X(_05751_));
 sky130_fd_sc_hd__nor2_4 _11114_ (.A(\CPU_Dmem_value_a5[11][9] ),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a211o_4 _11115_ (.A1(_05322_),
    .A2(_05748_),
    .B1(_05741_),
    .C1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__inv_2 _11116_ (.A(_05753_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_4 _11117_ (.A(\CPU_Dmem_value_a5[11][8] ),
    .B(_05751_),
    .Y(_05754_));
 sky130_fd_sc_hd__a211o_4 _11118_ (.A1(_05325_),
    .A2(_05748_),
    .B1(_05741_),
    .C1(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__inv_2 _11119_ (.A(_05755_),
    .Y(_01174_));
 sky130_fd_sc_hd__buf_2 _11120_ (.A(_05740_),
    .X(_05756_));
 sky130_fd_sc_hd__nor2_4 _11121_ (.A(\CPU_Dmem_value_a5[11][7] ),
    .B(_05751_),
    .Y(_05757_));
 sky130_fd_sc_hd__a211o_4 _11122_ (.A1(_05328_),
    .A2(_05748_),
    .B1(_05756_),
    .C1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__inv_2 _11123_ (.A(_05758_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_4 _11124_ (.A(\CPU_Dmem_value_a5[11][6] ),
    .B(_05751_),
    .Y(_05759_));
 sky130_fd_sc_hd__a211o_4 _11125_ (.A1(_05333_),
    .A2(_05748_),
    .B1(_05756_),
    .C1(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__inv_2 _11126_ (.A(_05760_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor2_4 _11127_ (.A(\CPU_Dmem_value_a5[11][5] ),
    .B(_05751_),
    .Y(_05761_));
 sky130_fd_sc_hd__a211o_4 _11128_ (.A1(_05336_),
    .A2(_05748_),
    .B1(_05756_),
    .C1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__inv_2 _11129_ (.A(_05762_),
    .Y(_01171_));
 sky130_fd_sc_hd__nor2_4 _11130_ (.A(\CPU_Dmem_value_a5[11][4] ),
    .B(_05751_),
    .Y(_05763_));
 sky130_fd_sc_hd__a211o_4 _11131_ (.A1(_05339_),
    .A2(_05695_),
    .B1(_05756_),
    .C1(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__inv_2 _11132_ (.A(_05764_),
    .Y(_01170_));
 sky130_fd_sc_hd__and2_4 _11133_ (.A(\CPU_Dmem_value_a5[11][3] ),
    .B(_05690_),
    .X(_05765_));
 sky130_fd_sc_hd__a211o_4 _11134_ (.A1(_05510_),
    .A2(_05693_),
    .B1(_05511_),
    .C1(_05765_),
    .X(_01169_));
 sky130_fd_sc_hd__nor2_4 _11135_ (.A(\CPU_Dmem_value_a5[11][2] ),
    .B(_05692_),
    .Y(_05766_));
 sky130_fd_sc_hd__a211o_4 _11136_ (.A1(_04787_),
    .A2(_05695_),
    .B1(_05756_),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__inv_2 _11137_ (.A(_05767_),
    .Y(_01168_));
 sky130_fd_sc_hd__buf_2 _11138_ (.A(_04888_),
    .X(_05768_));
 sky130_fd_sc_hd__and2_4 _11139_ (.A(\CPU_Dmem_value_a5[11][1] ),
    .B(_05690_),
    .X(_05769_));
 sky130_fd_sc_hd__a211o_4 _11140_ (.A1(_04976_),
    .A2(_05693_),
    .B1(_05768_),
    .C1(_05769_),
    .X(_01167_));
 sky130_fd_sc_hd__and2_4 _11141_ (.A(\CPU_Dmem_value_a5[11][0] ),
    .B(_05690_),
    .X(_05770_));
 sky130_fd_sc_hd__a211o_4 _11142_ (.A1(_04887_),
    .A2(_05693_),
    .B1(_05768_),
    .C1(_05770_),
    .X(_01166_));
 sky130_fd_sc_hd__or4_4 _11143_ (.A(_04650_),
    .B(_04651_),
    .C(_05605_),
    .D(_05067_),
    .X(_05771_));
 sky130_fd_sc_hd__buf_2 _11144_ (.A(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__nor2_4 _11145_ (.A(_05351_),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__buf_2 _11146_ (.A(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__buf_2 _11147_ (.A(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__buf_2 _11148_ (.A(_05774_),
    .X(_05776_));
 sky130_fd_sc_hd__nor2_4 _11149_ (.A(\CPU_Dmem_value_a5[12][31] ),
    .B(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__a211o_4 _11150_ (.A1(_05350_),
    .A2(_05775_),
    .B1(_05756_),
    .C1(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__inv_2 _11151_ (.A(_05778_),
    .Y(_01165_));
 sky130_fd_sc_hd__buf_2 _11152_ (.A(_05740_),
    .X(_05779_));
 sky130_fd_sc_hd__nor2_4 _11153_ (.A(\CPU_Dmem_value_a5[12][30] ),
    .B(_05776_),
    .Y(_05780_));
 sky130_fd_sc_hd__a211o_4 _11154_ (.A1(_04646_),
    .A2(_05775_),
    .B1(_05779_),
    .C1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__inv_2 _11155_ (.A(_05781_),
    .Y(_01164_));
 sky130_fd_sc_hd__buf_2 _11156_ (.A(_05773_),
    .X(_05782_));
 sky130_fd_sc_hd__buf_2 _11157_ (.A(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__buf_2 _11158_ (.A(_05774_),
    .X(_05784_));
 sky130_fd_sc_hd__nor2_4 _11159_ (.A(\CPU_Dmem_value_a5[12][29] ),
    .B(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__a211o_4 _11160_ (.A1(_04667_),
    .A2(_05783_),
    .B1(_05779_),
    .C1(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__inv_2 _11161_ (.A(_05786_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_4 _11162_ (.A(\CPU_Dmem_value_a5[12][28] ),
    .B(_05784_),
    .Y(_05787_));
 sky130_fd_sc_hd__a211o_4 _11163_ (.A1(_04671_),
    .A2(_05783_),
    .B1(_05779_),
    .C1(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__inv_2 _11164_ (.A(_05788_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_4 _11165_ (.A(\CPU_Dmem_value_a5[12][27] ),
    .B(_05784_),
    .Y(_05789_));
 sky130_fd_sc_hd__a211o_4 _11166_ (.A1(_04675_),
    .A2(_05783_),
    .B1(_05779_),
    .C1(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__inv_2 _11167_ (.A(_05790_),
    .Y(_01161_));
 sky130_fd_sc_hd__nor2_4 _11168_ (.A(\CPU_Dmem_value_a5[12][26] ),
    .B(_05784_),
    .Y(_05791_));
 sky130_fd_sc_hd__a211o_4 _11169_ (.A1(_04679_),
    .A2(_05783_),
    .B1(_05779_),
    .C1(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__inv_2 _11170_ (.A(_05792_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_4 _11171_ (.A(\CPU_Dmem_value_a5[12][25] ),
    .B(_05784_),
    .Y(_05793_));
 sky130_fd_sc_hd__a211o_4 _11172_ (.A1(_04685_),
    .A2(_05783_),
    .B1(_05779_),
    .C1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__inv_2 _11173_ (.A(_05794_),
    .Y(_01159_));
 sky130_fd_sc_hd__buf_2 _11174_ (.A(_05740_),
    .X(_05795_));
 sky130_fd_sc_hd__nor2_4 _11175_ (.A(\CPU_Dmem_value_a5[12][24] ),
    .B(_05784_),
    .Y(_05796_));
 sky130_fd_sc_hd__a211o_4 _11176_ (.A1(_04689_),
    .A2(_05783_),
    .B1(_05795_),
    .C1(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__inv_2 _11177_ (.A(_05797_),
    .Y(_01158_));
 sky130_fd_sc_hd__buf_2 _11178_ (.A(_05782_),
    .X(_05798_));
 sky130_fd_sc_hd__buf_2 _11179_ (.A(_05774_),
    .X(_05799_));
 sky130_fd_sc_hd__nor2_4 _11180_ (.A(\CPU_Dmem_value_a5[12][23] ),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__a211o_4 _11181_ (.A1(_04694_),
    .A2(_05798_),
    .B1(_05795_),
    .C1(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__inv_2 _11182_ (.A(_05801_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_4 _11183_ (.A(\CPU_Dmem_value_a5[12][22] ),
    .B(_05799_),
    .Y(_05802_));
 sky130_fd_sc_hd__a211o_4 _11184_ (.A1(_04698_),
    .A2(_05798_),
    .B1(_05795_),
    .C1(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__inv_2 _11185_ (.A(_05803_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_4 _11186_ (.A(\CPU_Dmem_value_a5[12][21] ),
    .B(_05799_),
    .Y(_05804_));
 sky130_fd_sc_hd__a211o_4 _11187_ (.A1(_04702_),
    .A2(_05798_),
    .B1(_05795_),
    .C1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__inv_2 _11188_ (.A(_05805_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_4 _11189_ (.A(\CPU_Dmem_value_a5[12][20] ),
    .B(_05799_),
    .Y(_05806_));
 sky130_fd_sc_hd__a211o_4 _11190_ (.A1(_04706_),
    .A2(_05798_),
    .B1(_05795_),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__inv_2 _11191_ (.A(_05807_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_4 _11192_ (.A(\CPU_Dmem_value_a5[12][19] ),
    .B(_05799_),
    .Y(_05808_));
 sky130_fd_sc_hd__a211o_4 _11193_ (.A1(_04712_),
    .A2(_05798_),
    .B1(_05795_),
    .C1(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__inv_2 _11194_ (.A(_05809_),
    .Y(_01153_));
 sky130_fd_sc_hd__buf_2 _11195_ (.A(_05740_),
    .X(_05810_));
 sky130_fd_sc_hd__nor2_4 _11196_ (.A(\CPU_Dmem_value_a5[12][18] ),
    .B(_05799_),
    .Y(_05811_));
 sky130_fd_sc_hd__a211o_4 _11197_ (.A1(_04716_),
    .A2(_05798_),
    .B1(_05810_),
    .C1(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__inv_2 _11198_ (.A(_05812_),
    .Y(_01152_));
 sky130_fd_sc_hd__buf_2 _11199_ (.A(_05774_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_2 _11200_ (.A(_05773_),
    .X(_05814_));
 sky130_fd_sc_hd__nor2_4 _11201_ (.A(\CPU_Dmem_value_a5[12][17] ),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__a211o_4 _11202_ (.A1(_04721_),
    .A2(_05813_),
    .B1(_05810_),
    .C1(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__inv_2 _11203_ (.A(_05816_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_4 _11204_ (.A(\CPU_Dmem_value_a5[12][16] ),
    .B(_05814_),
    .Y(_05817_));
 sky130_fd_sc_hd__a211o_4 _11205_ (.A1(_04725_),
    .A2(_05813_),
    .B1(_05810_),
    .C1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__inv_2 _11206_ (.A(_05818_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_4 _11207_ (.A(\CPU_Dmem_value_a5[12][15] ),
    .B(_05814_),
    .Y(_05819_));
 sky130_fd_sc_hd__a211o_4 _11208_ (.A1(_04729_),
    .A2(_05813_),
    .B1(_05810_),
    .C1(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__inv_2 _11209_ (.A(_05820_),
    .Y(_01149_));
 sky130_fd_sc_hd__nor2_4 _11210_ (.A(\CPU_Dmem_value_a5[12][14] ),
    .B(_05814_),
    .Y(_05821_));
 sky130_fd_sc_hd__a211o_4 _11211_ (.A1(_04733_),
    .A2(_05813_),
    .B1(_05810_),
    .C1(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__inv_2 _11212_ (.A(_05822_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_4 _11213_ (.A(\CPU_Dmem_value_a5[12][13] ),
    .B(_05814_),
    .Y(_05823_));
 sky130_fd_sc_hd__a211o_4 _11214_ (.A1(_04739_),
    .A2(_05813_),
    .B1(_05810_),
    .C1(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__inv_2 _11215_ (.A(_05824_),
    .Y(_01147_));
 sky130_fd_sc_hd__buf_2 _11216_ (.A(_05740_),
    .X(_05825_));
 sky130_fd_sc_hd__nor2_4 _11217_ (.A(\CPU_Dmem_value_a5[12][12] ),
    .B(_05814_),
    .Y(_05826_));
 sky130_fd_sc_hd__a211o_4 _11218_ (.A1(_04743_),
    .A2(_05813_),
    .B1(_05825_),
    .C1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__inv_2 _11219_ (.A(_05827_),
    .Y(_01146_));
 sky130_fd_sc_hd__buf_2 _11220_ (.A(_05774_),
    .X(_05828_));
 sky130_fd_sc_hd__buf_2 _11221_ (.A(_05773_),
    .X(_05829_));
 sky130_fd_sc_hd__nor2_4 _11222_ (.A(\CPU_Dmem_value_a5[12][11] ),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a211o_4 _11223_ (.A1(_04748_),
    .A2(_05828_),
    .B1(_05825_),
    .C1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__inv_2 _11224_ (.A(_05831_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_4 _11225_ (.A(\CPU_Dmem_value_a5[12][10] ),
    .B(_05829_),
    .Y(_05832_));
 sky130_fd_sc_hd__a211o_4 _11226_ (.A1(_04752_),
    .A2(_05828_),
    .B1(_05825_),
    .C1(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__inv_2 _11227_ (.A(_05833_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_4 _11228_ (.A(\CPU_Dmem_value_a5[12][9] ),
    .B(_05829_),
    .Y(_05834_));
 sky130_fd_sc_hd__a211o_4 _11229_ (.A1(_04756_),
    .A2(_05828_),
    .B1(_05825_),
    .C1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__inv_2 _11230_ (.A(_05835_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_4 _11231_ (.A(\CPU_Dmem_value_a5[12][8] ),
    .B(_05829_),
    .Y(_05836_));
 sky130_fd_sc_hd__a211o_4 _11232_ (.A1(_04760_),
    .A2(_05828_),
    .B1(_05825_),
    .C1(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__inv_2 _11233_ (.A(_05837_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_4 _11234_ (.A(\CPU_Dmem_value_a5[12][7] ),
    .B(_05829_),
    .Y(_05838_));
 sky130_fd_sc_hd__a211o_4 _11235_ (.A1(_04766_),
    .A2(_05828_),
    .B1(_05825_),
    .C1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__inv_2 _11236_ (.A(_05839_),
    .Y(_01141_));
 sky130_fd_sc_hd__buf_2 _11237_ (.A(_04659_),
    .X(_05840_));
 sky130_fd_sc_hd__buf_2 _11238_ (.A(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__nor2_4 _11239_ (.A(\CPU_Dmem_value_a5[12][6] ),
    .B(_05829_),
    .Y(_05842_));
 sky130_fd_sc_hd__a211o_4 _11240_ (.A1(_04770_),
    .A2(_05828_),
    .B1(_05841_),
    .C1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__inv_2 _11241_ (.A(_05843_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_4 _11242_ (.A(\CPU_Dmem_value_a5[12][5] ),
    .B(_05782_),
    .Y(_05844_));
 sky130_fd_sc_hd__a211o_4 _11243_ (.A1(_04775_),
    .A2(_05776_),
    .B1(_05841_),
    .C1(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__inv_2 _11244_ (.A(_05845_),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_4 _11245_ (.A(\CPU_Dmem_value_a5[12][4] ),
    .B(_05782_),
    .Y(_05846_));
 sky130_fd_sc_hd__a211o_4 _11246_ (.A1(_04779_),
    .A2(_05776_),
    .B1(_05841_),
    .C1(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__inv_2 _11247_ (.A(_05847_),
    .Y(_01138_));
 sky130_fd_sc_hd__inv_2 _11248_ (.A(\CPU_Dmem_value_a5[12][3] ),
    .Y(_05848_));
 sky130_fd_sc_hd__nor2_4 _11249_ (.A(_05848_),
    .B(_05775_),
    .Y(_05849_));
 sky130_fd_sc_hd__a211o_4 _11250_ (.A1(_05510_),
    .A2(_05775_),
    .B1(_05768_),
    .C1(_05849_),
    .X(_01137_));
 sky130_fd_sc_hd__inv_2 _11251_ (.A(\CPU_Dmem_value_a5[12][2] ),
    .Y(_05850_));
 sky130_fd_sc_hd__nor2_4 _11252_ (.A(_05850_),
    .B(_05775_),
    .Y(_05851_));
 sky130_fd_sc_hd__a211o_4 _11253_ (.A1(_05147_),
    .A2(_05775_),
    .B1(_05768_),
    .C1(_05851_),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_4 _11254_ (.A(\CPU_Dmem_value_a5[12][1] ),
    .B(_05782_),
    .Y(_05852_));
 sky130_fd_sc_hd__a211o_4 _11255_ (.A1(_04793_),
    .A2(_05776_),
    .B1(_05841_),
    .C1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__inv_2 _11256_ (.A(_05853_),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_4 _11257_ (.A(\CPU_Dmem_value_a5[12][0] ),
    .B(_05782_),
    .Y(_05854_));
 sky130_fd_sc_hd__a211o_4 _11258_ (.A1(_04797_),
    .A2(_05776_),
    .B1(_05841_),
    .C1(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__inv_2 _11259_ (.A(_05855_),
    .Y(_01134_));
 sky130_fd_sc_hd__or4_4 _11260_ (.A(_04650_),
    .B(_04804_),
    .C(_05605_),
    .D(_05067_),
    .X(_05856_));
 sky130_fd_sc_hd__or2_4 _11261_ (.A(_05351_),
    .B(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__inv_2 _11262_ (.A(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__buf_2 _11263_ (.A(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__buf_2 _11264_ (.A(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__buf_2 _11265_ (.A(_05858_),
    .X(_05861_));
 sky130_fd_sc_hd__nor2_4 _11266_ (.A(\CPU_Dmem_value_a5[13][31] ),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__a211o_4 _11267_ (.A1(_04801_),
    .A2(_05860_),
    .B1(_05841_),
    .C1(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__inv_2 _11268_ (.A(_05863_),
    .Y(_01133_));
 sky130_fd_sc_hd__buf_2 _11269_ (.A(_05840_),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_4 _11270_ (.A(\CPU_Dmem_value_a5[13][30] ),
    .B(_05861_),
    .Y(_05865_));
 sky130_fd_sc_hd__a211o_4 _11271_ (.A1(_04646_),
    .A2(_05860_),
    .B1(_05864_),
    .C1(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__inv_2 _11272_ (.A(_05866_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_4 _11273_ (.A(\CPU_Dmem_value_a5[13][29] ),
    .B(_05861_),
    .Y(_05867_));
 sky130_fd_sc_hd__a211o_4 _11274_ (.A1(_04667_),
    .A2(_05860_),
    .B1(_05864_),
    .C1(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__inv_2 _11275_ (.A(_05868_),
    .Y(_01131_));
 sky130_fd_sc_hd__buf_2 _11276_ (.A(_05859_),
    .X(_05869_));
 sky130_fd_sc_hd__nor2_4 _11277_ (.A(\CPU_Dmem_value_a5[13][28] ),
    .B(_05861_),
    .Y(_05870_));
 sky130_fd_sc_hd__a211o_4 _11278_ (.A1(_04671_),
    .A2(_05869_),
    .B1(_05864_),
    .C1(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__inv_2 _11279_ (.A(_05871_),
    .Y(_01130_));
 sky130_fd_sc_hd__buf_2 _11280_ (.A(_05858_),
    .X(_05872_));
 sky130_fd_sc_hd__nor2_4 _11281_ (.A(\CPU_Dmem_value_a5[13][27] ),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__a211o_4 _11282_ (.A1(_04675_),
    .A2(_05869_),
    .B1(_05864_),
    .C1(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__inv_2 _11283_ (.A(_05874_),
    .Y(_01129_));
 sky130_fd_sc_hd__nor2_4 _11284_ (.A(\CPU_Dmem_value_a5[13][26] ),
    .B(_05872_),
    .Y(_05875_));
 sky130_fd_sc_hd__a211o_4 _11285_ (.A1(_04679_),
    .A2(_05869_),
    .B1(_05864_),
    .C1(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__inv_2 _11286_ (.A(_05876_),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_4 _11287_ (.A(\CPU_Dmem_value_a5[13][25] ),
    .B(_05872_),
    .Y(_05877_));
 sky130_fd_sc_hd__a211o_4 _11288_ (.A1(_04685_),
    .A2(_05869_),
    .B1(_05864_),
    .C1(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__inv_2 _11289_ (.A(_05878_),
    .Y(_01127_));
 sky130_fd_sc_hd__buf_2 _11290_ (.A(_05840_),
    .X(_05879_));
 sky130_fd_sc_hd__nor2_4 _11291_ (.A(\CPU_Dmem_value_a5[13][24] ),
    .B(_05872_),
    .Y(_05880_));
 sky130_fd_sc_hd__a211o_4 _11292_ (.A1(_04689_),
    .A2(_05869_),
    .B1(_05879_),
    .C1(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__inv_2 _11293_ (.A(_05881_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_4 _11294_ (.A(\CPU_Dmem_value_a5[13][23] ),
    .B(_05872_),
    .Y(_05882_));
 sky130_fd_sc_hd__a211o_4 _11295_ (.A1(_04694_),
    .A2(_05869_),
    .B1(_05879_),
    .C1(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__inv_2 _11296_ (.A(_05883_),
    .Y(_01125_));
 sky130_fd_sc_hd__buf_2 _11297_ (.A(_05859_),
    .X(_05884_));
 sky130_fd_sc_hd__nor2_4 _11298_ (.A(\CPU_Dmem_value_a5[13][22] ),
    .B(_05872_),
    .Y(_05885_));
 sky130_fd_sc_hd__a211o_4 _11299_ (.A1(_04698_),
    .A2(_05884_),
    .B1(_05879_),
    .C1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__inv_2 _11300_ (.A(_05886_),
    .Y(_01124_));
 sky130_fd_sc_hd__buf_2 _11301_ (.A(_05858_),
    .X(_05887_));
 sky130_fd_sc_hd__nor2_4 _11302_ (.A(\CPU_Dmem_value_a5[13][21] ),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__a211o_4 _11303_ (.A1(_04702_),
    .A2(_05884_),
    .B1(_05879_),
    .C1(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__inv_2 _11304_ (.A(_05889_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_4 _11305_ (.A(\CPU_Dmem_value_a5[13][20] ),
    .B(_05887_),
    .Y(_05890_));
 sky130_fd_sc_hd__a211o_4 _11306_ (.A1(_04706_),
    .A2(_05884_),
    .B1(_05879_),
    .C1(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__inv_2 _11307_ (.A(_05891_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_4 _11308_ (.A(\CPU_Dmem_value_a5[13][19] ),
    .B(_05887_),
    .Y(_05892_));
 sky130_fd_sc_hd__a211o_4 _11309_ (.A1(_04712_),
    .A2(_05884_),
    .B1(_05879_),
    .C1(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__inv_2 _11310_ (.A(_05893_),
    .Y(_01121_));
 sky130_fd_sc_hd__buf_2 _11311_ (.A(_05840_),
    .X(_05894_));
 sky130_fd_sc_hd__nor2_4 _11312_ (.A(\CPU_Dmem_value_a5[13][18] ),
    .B(_05887_),
    .Y(_05895_));
 sky130_fd_sc_hd__a211o_4 _11313_ (.A1(_04716_),
    .A2(_05884_),
    .B1(_05894_),
    .C1(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__inv_2 _11314_ (.A(_05896_),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_4 _11315_ (.A(\CPU_Dmem_value_a5[13][17] ),
    .B(_05887_),
    .Y(_05897_));
 sky130_fd_sc_hd__a211o_4 _11316_ (.A1(_04721_),
    .A2(_05884_),
    .B1(_05894_),
    .C1(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__inv_2 _11317_ (.A(_05898_),
    .Y(_01119_));
 sky130_fd_sc_hd__buf_2 _11318_ (.A(_05859_),
    .X(_05899_));
 sky130_fd_sc_hd__nor2_4 _11319_ (.A(\CPU_Dmem_value_a5[13][16] ),
    .B(_05887_),
    .Y(_05900_));
 sky130_fd_sc_hd__a211o_4 _11320_ (.A1(_04725_),
    .A2(_05899_),
    .B1(_05894_),
    .C1(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__inv_2 _11321_ (.A(_05901_),
    .Y(_01118_));
 sky130_fd_sc_hd__buf_2 _11322_ (.A(_05858_),
    .X(_05902_));
 sky130_fd_sc_hd__nor2_4 _11323_ (.A(\CPU_Dmem_value_a5[13][15] ),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__a211o_4 _11324_ (.A1(_04729_),
    .A2(_05899_),
    .B1(_05894_),
    .C1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__inv_2 _11325_ (.A(_05904_),
    .Y(_01117_));
 sky130_fd_sc_hd__nor2_4 _11326_ (.A(\CPU_Dmem_value_a5[13][14] ),
    .B(_05902_),
    .Y(_05905_));
 sky130_fd_sc_hd__a211o_4 _11327_ (.A1(_04733_),
    .A2(_05899_),
    .B1(_05894_),
    .C1(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__inv_2 _11328_ (.A(_05906_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_4 _11329_ (.A(\CPU_Dmem_value_a5[13][13] ),
    .B(_05902_),
    .Y(_05907_));
 sky130_fd_sc_hd__a211o_4 _11330_ (.A1(_04739_),
    .A2(_05899_),
    .B1(_05894_),
    .C1(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__inv_2 _11331_ (.A(_05908_),
    .Y(_01115_));
 sky130_fd_sc_hd__buf_2 _11332_ (.A(_05840_),
    .X(_05909_));
 sky130_fd_sc_hd__nor2_4 _11333_ (.A(\CPU_Dmem_value_a5[13][12] ),
    .B(_05902_),
    .Y(_05910_));
 sky130_fd_sc_hd__a211o_4 _11334_ (.A1(_04743_),
    .A2(_05899_),
    .B1(_05909_),
    .C1(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__inv_2 _11335_ (.A(_05911_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_4 _11336_ (.A(\CPU_Dmem_value_a5[13][11] ),
    .B(_05902_),
    .Y(_05912_));
 sky130_fd_sc_hd__a211o_4 _11337_ (.A1(_04748_),
    .A2(_05899_),
    .B1(_05909_),
    .C1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__inv_2 _11338_ (.A(_05913_),
    .Y(_01113_));
 sky130_fd_sc_hd__buf_2 _11339_ (.A(_05859_),
    .X(_05914_));
 sky130_fd_sc_hd__nor2_4 _11340_ (.A(\CPU_Dmem_value_a5[13][10] ),
    .B(_05902_),
    .Y(_05915_));
 sky130_fd_sc_hd__a211o_4 _11341_ (.A1(_04752_),
    .A2(_05914_),
    .B1(_05909_),
    .C1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__inv_2 _11342_ (.A(_05916_),
    .Y(_01112_));
 sky130_fd_sc_hd__buf_2 _11343_ (.A(_05858_),
    .X(_05917_));
 sky130_fd_sc_hd__nor2_4 _11344_ (.A(\CPU_Dmem_value_a5[13][9] ),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a211o_4 _11345_ (.A1(_04756_),
    .A2(_05914_),
    .B1(_05909_),
    .C1(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__inv_2 _11346_ (.A(_05919_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_4 _11347_ (.A(\CPU_Dmem_value_a5[13][8] ),
    .B(_05917_),
    .Y(_05920_));
 sky130_fd_sc_hd__a211o_4 _11348_ (.A1(_04760_),
    .A2(_05914_),
    .B1(_05909_),
    .C1(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__inv_2 _11349_ (.A(_05921_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_4 _11350_ (.A(\CPU_Dmem_value_a5[13][7] ),
    .B(_05917_),
    .Y(_05922_));
 sky130_fd_sc_hd__a211o_4 _11351_ (.A1(_04766_),
    .A2(_05914_),
    .B1(_05909_),
    .C1(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__inv_2 _11352_ (.A(_05923_),
    .Y(_01109_));
 sky130_fd_sc_hd__buf_2 _11353_ (.A(_05840_),
    .X(_05924_));
 sky130_fd_sc_hd__nor2_4 _11354_ (.A(\CPU_Dmem_value_a5[13][6] ),
    .B(_05917_),
    .Y(_05925_));
 sky130_fd_sc_hd__a211o_4 _11355_ (.A1(_04770_),
    .A2(_05914_),
    .B1(_05924_),
    .C1(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__inv_2 _11356_ (.A(_05926_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_4 _11357_ (.A(\CPU_Dmem_value_a5[13][5] ),
    .B(_05917_),
    .Y(_05927_));
 sky130_fd_sc_hd__a211o_4 _11358_ (.A1(_04775_),
    .A2(_05914_),
    .B1(_05924_),
    .C1(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__inv_2 _11359_ (.A(_05928_),
    .Y(_01107_));
 sky130_fd_sc_hd__nor2_4 _11360_ (.A(\CPU_Dmem_value_a5[13][4] ),
    .B(_05917_),
    .Y(_05929_));
 sky130_fd_sc_hd__a211o_4 _11361_ (.A1(_04779_),
    .A2(_05861_),
    .B1(_05924_),
    .C1(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__inv_2 _11362_ (.A(_05930_),
    .Y(_01106_));
 sky130_fd_sc_hd__and2_4 _11363_ (.A(\CPU_Dmem_value_a5[13][3] ),
    .B(_05857_),
    .X(_05931_));
 sky130_fd_sc_hd__a211o_4 _11364_ (.A1(_05510_),
    .A2(_05860_),
    .B1(_05768_),
    .C1(_05931_),
    .X(_01105_));
 sky130_fd_sc_hd__and2_4 _11365_ (.A(\CPU_Dmem_value_a5[13][2] ),
    .B(_05857_),
    .X(_05932_));
 sky130_fd_sc_hd__a211o_4 _11366_ (.A1(_05147_),
    .A2(_05860_),
    .B1(_05768_),
    .C1(_05932_),
    .X(_01104_));
 sky130_fd_sc_hd__nor2_4 _11367_ (.A(\CPU_Dmem_value_a5[13][1] ),
    .B(_05859_),
    .Y(_05933_));
 sky130_fd_sc_hd__a211o_4 _11368_ (.A1(_04793_),
    .A2(_05861_),
    .B1(_05924_),
    .C1(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__inv_2 _11369_ (.A(_05934_),
    .Y(_01103_));
 sky130_fd_sc_hd__buf_2 _11370_ (.A(_04661_),
    .X(_05935_));
 sky130_fd_sc_hd__and2_4 _11371_ (.A(\CPU_Dmem_value_a5[13][0] ),
    .B(_05857_),
    .X(_05936_));
 sky130_fd_sc_hd__a211o_4 _11372_ (.A1(\CPU_dmem_wr_data_a4[0] ),
    .A2(_05860_),
    .B1(_05935_),
    .C1(_05936_),
    .X(_01102_));
 sky130_fd_sc_hd__or4_4 _11373_ (.A(_04893_),
    .B(_04651_),
    .C(_05605_),
    .D(_05067_),
    .X(_05937_));
 sky130_fd_sc_hd__buf_2 _11374_ (.A(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__nor2_4 _11375_ (.A(_05351_),
    .B(_05938_),
    .Y(_05939_));
 sky130_fd_sc_hd__buf_2 _11376_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__buf_2 _11377_ (.A(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__buf_2 _11378_ (.A(_05939_),
    .X(_05942_));
 sky130_fd_sc_hd__buf_2 _11379_ (.A(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__nor2_4 _11380_ (.A(\CPU_Dmem_value_a5[14][31] ),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__a211o_4 _11381_ (.A1(_04801_),
    .A2(_05941_),
    .B1(_05924_),
    .C1(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__inv_2 _11382_ (.A(_05945_),
    .Y(_01101_));
 sky130_fd_sc_hd__buf_2 _11383_ (.A(_05942_),
    .X(_05946_));
 sky130_fd_sc_hd__nor2_4 _11384_ (.A(\CPU_Dmem_value_a5[14][30] ),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__a211o_4 _11385_ (.A1(_04646_),
    .A2(_05941_),
    .B1(_05924_),
    .C1(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__inv_2 _11386_ (.A(_05948_),
    .Y(_01100_));
 sky130_fd_sc_hd__buf_2 _11387_ (.A(_04659_),
    .X(_05949_));
 sky130_fd_sc_hd__buf_2 _11388_ (.A(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_4 _11389_ (.A(\CPU_Dmem_value_a5[14][29] ),
    .B(_05946_),
    .Y(_05951_));
 sky130_fd_sc_hd__a211o_4 _11390_ (.A1(_04667_),
    .A2(_05941_),
    .B1(_05950_),
    .C1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__inv_2 _11391_ (.A(_05952_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_4 _11392_ (.A(\CPU_Dmem_value_a5[14][28] ),
    .B(_05946_),
    .Y(_05953_));
 sky130_fd_sc_hd__a211o_4 _11393_ (.A1(_04671_),
    .A2(_05941_),
    .B1(_05950_),
    .C1(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__inv_2 _11394_ (.A(_05954_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_4 _11395_ (.A(\CPU_Dmem_value_a5[14][27] ),
    .B(_05946_),
    .Y(_05955_));
 sky130_fd_sc_hd__a211o_4 _11396_ (.A1(_04675_),
    .A2(_05941_),
    .B1(_05950_),
    .C1(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__inv_2 _11397_ (.A(_05956_),
    .Y(_01097_));
 sky130_fd_sc_hd__nor2_4 _11398_ (.A(\CPU_Dmem_value_a5[14][26] ),
    .B(_05946_),
    .Y(_05957_));
 sky130_fd_sc_hd__a211o_4 _11399_ (.A1(_04679_),
    .A2(_05941_),
    .B1(_05950_),
    .C1(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__inv_2 _11400_ (.A(_05958_),
    .Y(_01096_));
 sky130_fd_sc_hd__buf_2 _11401_ (.A(_05942_),
    .X(_05959_));
 sky130_fd_sc_hd__nor2_4 _11402_ (.A(\CPU_Dmem_value_a5[14][25] ),
    .B(_05946_),
    .Y(_05960_));
 sky130_fd_sc_hd__a211o_4 _11403_ (.A1(_04685_),
    .A2(_05959_),
    .B1(_05950_),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__inv_2 _11404_ (.A(_05961_),
    .Y(_01095_));
 sky130_fd_sc_hd__buf_2 _11405_ (.A(_05942_),
    .X(_05962_));
 sky130_fd_sc_hd__nor2_4 _11406_ (.A(\CPU_Dmem_value_a5[14][24] ),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a211o_4 _11407_ (.A1(_04689_),
    .A2(_05959_),
    .B1(_05950_),
    .C1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__inv_2 _11408_ (.A(_05964_),
    .Y(_01094_));
 sky130_fd_sc_hd__buf_2 _11409_ (.A(_05949_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_4 _11410_ (.A(\CPU_Dmem_value_a5[14][23] ),
    .B(_05962_),
    .Y(_05966_));
 sky130_fd_sc_hd__a211o_4 _11411_ (.A1(_04694_),
    .A2(_05959_),
    .B1(_05965_),
    .C1(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__inv_2 _11412_ (.A(_05967_),
    .Y(_01093_));
 sky130_fd_sc_hd__nor2_4 _11413_ (.A(\CPU_Dmem_value_a5[14][22] ),
    .B(_05962_),
    .Y(_05968_));
 sky130_fd_sc_hd__a211o_4 _11414_ (.A1(_04698_),
    .A2(_05959_),
    .B1(_05965_),
    .C1(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__inv_2 _11415_ (.A(_05969_),
    .Y(_01092_));
 sky130_fd_sc_hd__nor2_4 _11416_ (.A(\CPU_Dmem_value_a5[14][21] ),
    .B(_05962_),
    .Y(_05970_));
 sky130_fd_sc_hd__a211o_4 _11417_ (.A1(_04702_),
    .A2(_05959_),
    .B1(_05965_),
    .C1(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__inv_2 _11418_ (.A(_05971_),
    .Y(_01091_));
 sky130_fd_sc_hd__nor2_4 _11419_ (.A(\CPU_Dmem_value_a5[14][20] ),
    .B(_05962_),
    .Y(_05972_));
 sky130_fd_sc_hd__a211o_4 _11420_ (.A1(_04706_),
    .A2(_05959_),
    .B1(_05965_),
    .C1(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__inv_2 _11421_ (.A(_05973_),
    .Y(_01090_));
 sky130_fd_sc_hd__buf_2 _11422_ (.A(_05942_),
    .X(_05974_));
 sky130_fd_sc_hd__nor2_4 _11423_ (.A(\CPU_Dmem_value_a5[14][19] ),
    .B(_05962_),
    .Y(_05975_));
 sky130_fd_sc_hd__a211o_4 _11424_ (.A1(_04712_),
    .A2(_05974_),
    .B1(_05965_),
    .C1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__inv_2 _11425_ (.A(_05976_),
    .Y(_01089_));
 sky130_fd_sc_hd__buf_2 _11426_ (.A(_05939_),
    .X(_05977_));
 sky130_fd_sc_hd__nor2_4 _11427_ (.A(\CPU_Dmem_value_a5[14][18] ),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__a211o_4 _11428_ (.A1(_04716_),
    .A2(_05974_),
    .B1(_05965_),
    .C1(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__inv_2 _11429_ (.A(_05979_),
    .Y(_01088_));
 sky130_fd_sc_hd__buf_2 _11430_ (.A(_05949_),
    .X(_05980_));
 sky130_fd_sc_hd__nor2_4 _11431_ (.A(\CPU_Dmem_value_a5[14][17] ),
    .B(_05977_),
    .Y(_05981_));
 sky130_fd_sc_hd__a211o_4 _11432_ (.A1(_04721_),
    .A2(_05974_),
    .B1(_05980_),
    .C1(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__inv_2 _11433_ (.A(_05982_),
    .Y(_01087_));
 sky130_fd_sc_hd__nor2_4 _11434_ (.A(\CPU_Dmem_value_a5[14][16] ),
    .B(_05977_),
    .Y(_05983_));
 sky130_fd_sc_hd__a211o_4 _11435_ (.A1(_04725_),
    .A2(_05974_),
    .B1(_05980_),
    .C1(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__inv_2 _11436_ (.A(_05984_),
    .Y(_01086_));
 sky130_fd_sc_hd__nor2_4 _11437_ (.A(\CPU_Dmem_value_a5[14][15] ),
    .B(_05977_),
    .Y(_05985_));
 sky130_fd_sc_hd__a211o_4 _11438_ (.A1(_04729_),
    .A2(_05974_),
    .B1(_05980_),
    .C1(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__inv_2 _11439_ (.A(_05986_),
    .Y(_01085_));
 sky130_fd_sc_hd__nor2_4 _11440_ (.A(\CPU_Dmem_value_a5[14][14] ),
    .B(_05977_),
    .Y(_05987_));
 sky130_fd_sc_hd__a211o_4 _11441_ (.A1(_04733_),
    .A2(_05974_),
    .B1(_05980_),
    .C1(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__inv_2 _11442_ (.A(_05988_),
    .Y(_01084_));
 sky130_fd_sc_hd__buf_2 _11443_ (.A(_05942_),
    .X(_05989_));
 sky130_fd_sc_hd__nor2_4 _11444_ (.A(\CPU_Dmem_value_a5[14][13] ),
    .B(_05977_),
    .Y(_05990_));
 sky130_fd_sc_hd__a211o_4 _11445_ (.A1(_04739_),
    .A2(_05989_),
    .B1(_05980_),
    .C1(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__inv_2 _11446_ (.A(_05991_),
    .Y(_01083_));
 sky130_fd_sc_hd__buf_2 _11447_ (.A(_05939_),
    .X(_05992_));
 sky130_fd_sc_hd__nor2_4 _11448_ (.A(\CPU_Dmem_value_a5[14][12] ),
    .B(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__a211o_4 _11449_ (.A1(_04743_),
    .A2(_05989_),
    .B1(_05980_),
    .C1(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__inv_2 _11450_ (.A(_05994_),
    .Y(_01082_));
 sky130_fd_sc_hd__buf_2 _11451_ (.A(_05949_),
    .X(_05995_));
 sky130_fd_sc_hd__nor2_4 _11452_ (.A(\CPU_Dmem_value_a5[14][11] ),
    .B(_05992_),
    .Y(_05996_));
 sky130_fd_sc_hd__a211o_4 _11453_ (.A1(_04748_),
    .A2(_05989_),
    .B1(_05995_),
    .C1(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__inv_2 _11454_ (.A(_05997_),
    .Y(_01081_));
 sky130_fd_sc_hd__nor2_4 _11455_ (.A(\CPU_Dmem_value_a5[14][10] ),
    .B(_05992_),
    .Y(_05998_));
 sky130_fd_sc_hd__a211o_4 _11456_ (.A1(_04752_),
    .A2(_05989_),
    .B1(_05995_),
    .C1(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__inv_2 _11457_ (.A(_05999_),
    .Y(_01080_));
 sky130_fd_sc_hd__nor2_4 _11458_ (.A(\CPU_Dmem_value_a5[14][9] ),
    .B(_05992_),
    .Y(_06000_));
 sky130_fd_sc_hd__a211o_4 _11459_ (.A1(_04756_),
    .A2(_05989_),
    .B1(_05995_),
    .C1(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__inv_2 _11460_ (.A(_06001_),
    .Y(_01079_));
 sky130_fd_sc_hd__nor2_4 _11461_ (.A(\CPU_Dmem_value_a5[14][8] ),
    .B(_05992_),
    .Y(_06002_));
 sky130_fd_sc_hd__a211o_4 _11462_ (.A1(_04760_),
    .A2(_05989_),
    .B1(_05995_),
    .C1(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__inv_2 _11463_ (.A(_06003_),
    .Y(_01078_));
 sky130_fd_sc_hd__nor2_4 _11464_ (.A(\CPU_Dmem_value_a5[14][7] ),
    .B(_05992_),
    .Y(_06004_));
 sky130_fd_sc_hd__a211o_4 _11465_ (.A1(_04766_),
    .A2(_05943_),
    .B1(_05995_),
    .C1(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__inv_2 _11466_ (.A(_06005_),
    .Y(_01077_));
 sky130_fd_sc_hd__nor2_4 _11467_ (.A(\CPU_Dmem_value_a5[14][6] ),
    .B(_05940_),
    .Y(_06006_));
 sky130_fd_sc_hd__a211o_4 _11468_ (.A1(_04770_),
    .A2(_05943_),
    .B1(_05995_),
    .C1(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__inv_2 _11469_ (.A(_06007_),
    .Y(_01076_));
 sky130_fd_sc_hd__buf_2 _11470_ (.A(_05949_),
    .X(_06008_));
 sky130_fd_sc_hd__nor2_4 _11471_ (.A(\CPU_Dmem_value_a5[14][5] ),
    .B(_05940_),
    .Y(_06009_));
 sky130_fd_sc_hd__a211o_4 _11472_ (.A1(_04775_),
    .A2(_05943_),
    .B1(_06008_),
    .C1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__inv_2 _11473_ (.A(_06010_),
    .Y(_01075_));
 sky130_fd_sc_hd__nor2_4 _11474_ (.A(\CPU_Dmem_value_a5[14][4] ),
    .B(_05940_),
    .Y(_06011_));
 sky130_fd_sc_hd__a211o_4 _11475_ (.A1(_04779_),
    .A2(_05943_),
    .B1(_06008_),
    .C1(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__inv_2 _11476_ (.A(_06012_),
    .Y(_01074_));
 sky130_fd_sc_hd__buf_2 _11477_ (.A(_05940_),
    .X(_06013_));
 sky130_fd_sc_hd__inv_2 _11478_ (.A(\CPU_Dmem_value_a5[14][3] ),
    .Y(_06014_));
 sky130_fd_sc_hd__nor2_4 _11479_ (.A(_06014_),
    .B(_06013_),
    .Y(_06015_));
 sky130_fd_sc_hd__a211o_4 _11480_ (.A1(\CPU_dmem_wr_data_a4[3] ),
    .A2(_06013_),
    .B1(_05935_),
    .C1(_06015_),
    .X(_01073_));
 sky130_fd_sc_hd__inv_2 _11481_ (.A(\CPU_Dmem_value_a5[14][2] ),
    .Y(_06016_));
 sky130_fd_sc_hd__nor2_4 _11482_ (.A(_06016_),
    .B(_06013_),
    .Y(_06017_));
 sky130_fd_sc_hd__a211o_4 _11483_ (.A1(\CPU_dmem_wr_data_a4[2] ),
    .A2(_06013_),
    .B1(_05935_),
    .C1(_06017_),
    .X(_01072_));
 sky130_fd_sc_hd__inv_2 _11484_ (.A(\CPU_Dmem_value_a5[14][1] ),
    .Y(_06018_));
 sky130_fd_sc_hd__nor2_4 _11485_ (.A(_06018_),
    .B(_06013_),
    .Y(_06019_));
 sky130_fd_sc_hd__a211o_4 _11486_ (.A1(\CPU_dmem_wr_data_a4[1] ),
    .A2(_06013_),
    .B1(_05935_),
    .C1(_06019_),
    .X(_01071_));
 sky130_fd_sc_hd__nor2_4 _11487_ (.A(\CPU_Dmem_value_a5[14][0] ),
    .B(_05940_),
    .Y(_06020_));
 sky130_fd_sc_hd__a211o_4 _11488_ (.A1(_04797_),
    .A2(_05943_),
    .B1(_06008_),
    .C1(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__inv_2 _11489_ (.A(_06021_),
    .Y(_01070_));
 sky130_fd_sc_hd__or4_4 _11490_ (.A(_04892_),
    .B(_04803_),
    .C(_05605_),
    .D(_05066_),
    .X(_06022_));
 sky130_fd_sc_hd__or2_4 _11491_ (.A(_04648_),
    .B(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__buf_2 _11493_ (.A(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__buf_2 _11494_ (.A(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__buf_2 _11495_ (.A(_06025_),
    .X(_06027_));
 sky130_fd_sc_hd__nor2_4 _11496_ (.A(\CPU_Dmem_value_a5[15][31] ),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a211o_4 _11497_ (.A1(_04801_),
    .A2(_06026_),
    .B1(_06008_),
    .C1(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__inv_2 _11498_ (.A(_06029_),
    .Y(_01069_));
 sky130_fd_sc_hd__nor2_4 _11499_ (.A(\CPU_Dmem_value_a5[15][30] ),
    .B(_06027_),
    .Y(_06030_));
 sky130_fd_sc_hd__a211o_4 _11500_ (.A1(_04646_),
    .A2(_06026_),
    .B1(_06008_),
    .C1(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__inv_2 _11501_ (.A(_06031_),
    .Y(_01068_));
 sky130_fd_sc_hd__buf_2 _11502_ (.A(_06025_),
    .X(_06032_));
 sky130_fd_sc_hd__nor2_4 _11503_ (.A(\CPU_Dmem_value_a5[15][29] ),
    .B(_06027_),
    .Y(_06033_));
 sky130_fd_sc_hd__a211o_4 _11504_ (.A1(_04667_),
    .A2(_06032_),
    .B1(_06008_),
    .C1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__inv_2 _11505_ (.A(_06034_),
    .Y(_01067_));
 sky130_fd_sc_hd__buf_2 _11506_ (.A(_05949_),
    .X(_06035_));
 sky130_fd_sc_hd__nor2_4 _11507_ (.A(\CPU_Dmem_value_a5[15][28] ),
    .B(_06027_),
    .Y(_06036_));
 sky130_fd_sc_hd__a211o_4 _11508_ (.A1(_04671_),
    .A2(_06032_),
    .B1(_06035_),
    .C1(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__inv_2 _11509_ (.A(_06037_),
    .Y(_01066_));
 sky130_fd_sc_hd__buf_2 _11510_ (.A(_06024_),
    .X(_06038_));
 sky130_fd_sc_hd__nor2_4 _11511_ (.A(\CPU_Dmem_value_a5[15][27] ),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__a211o_4 _11512_ (.A1(_04675_),
    .A2(_06032_),
    .B1(_06035_),
    .C1(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__inv_2 _11513_ (.A(_06040_),
    .Y(_01065_));
 sky130_fd_sc_hd__nor2_4 _11514_ (.A(\CPU_Dmem_value_a5[15][26] ),
    .B(_06038_),
    .Y(_06041_));
 sky130_fd_sc_hd__a211o_4 _11515_ (.A1(_04679_),
    .A2(_06032_),
    .B1(_06035_),
    .C1(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__inv_2 _11516_ (.A(_06042_),
    .Y(_01064_));
 sky130_fd_sc_hd__nor2_4 _11517_ (.A(\CPU_Dmem_value_a5[15][25] ),
    .B(_06038_),
    .Y(_06043_));
 sky130_fd_sc_hd__a211o_4 _11518_ (.A1(_04685_),
    .A2(_06032_),
    .B1(_06035_),
    .C1(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__inv_2 _11519_ (.A(_06044_),
    .Y(_01063_));
 sky130_fd_sc_hd__nor2_4 _11520_ (.A(\CPU_Dmem_value_a5[15][24] ),
    .B(_06038_),
    .Y(_06045_));
 sky130_fd_sc_hd__a211o_4 _11521_ (.A1(_04689_),
    .A2(_06032_),
    .B1(_06035_),
    .C1(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__inv_2 _11522_ (.A(_06046_),
    .Y(_01062_));
 sky130_fd_sc_hd__buf_2 _11523_ (.A(_06025_),
    .X(_06047_));
 sky130_fd_sc_hd__nor2_4 _11524_ (.A(\CPU_Dmem_value_a5[15][23] ),
    .B(_06038_),
    .Y(_06048_));
 sky130_fd_sc_hd__a211o_4 _11525_ (.A1(_04694_),
    .A2(_06047_),
    .B1(_06035_),
    .C1(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__inv_2 _11526_ (.A(_06049_),
    .Y(_01061_));
 sky130_fd_sc_hd__buf_2 _11527_ (.A(_04660_),
    .X(_06050_));
 sky130_fd_sc_hd__nor2_4 _11528_ (.A(\CPU_Dmem_value_a5[15][22] ),
    .B(_06038_),
    .Y(_06051_));
 sky130_fd_sc_hd__a211o_4 _11529_ (.A1(_04698_),
    .A2(_06047_),
    .B1(_06050_),
    .C1(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__inv_2 _11530_ (.A(_06052_),
    .Y(_01060_));
 sky130_fd_sc_hd__buf_2 _11531_ (.A(_06024_),
    .X(_06053_));
 sky130_fd_sc_hd__nor2_4 _11532_ (.A(\CPU_Dmem_value_a5[15][21] ),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a211o_4 _11533_ (.A1(_04702_),
    .A2(_06047_),
    .B1(_06050_),
    .C1(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__inv_2 _11534_ (.A(_06055_),
    .Y(_01059_));
 sky130_fd_sc_hd__nor2_4 _11535_ (.A(\CPU_Dmem_value_a5[15][20] ),
    .B(_06053_),
    .Y(_06056_));
 sky130_fd_sc_hd__a211o_4 _11536_ (.A1(_04706_),
    .A2(_06047_),
    .B1(_06050_),
    .C1(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__inv_2 _11537_ (.A(_06057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nor2_4 _11538_ (.A(\CPU_Dmem_value_a5[15][19] ),
    .B(_06053_),
    .Y(_06058_));
 sky130_fd_sc_hd__a211o_4 _11539_ (.A1(_04712_),
    .A2(_06047_),
    .B1(_06050_),
    .C1(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(_06059_),
    .Y(_01057_));
 sky130_fd_sc_hd__nor2_4 _11541_ (.A(\CPU_Dmem_value_a5[15][18] ),
    .B(_06053_),
    .Y(_06060_));
 sky130_fd_sc_hd__a211o_4 _11542_ (.A1(_04716_),
    .A2(_06047_),
    .B1(_06050_),
    .C1(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__inv_2 _11543_ (.A(_06061_),
    .Y(_01056_));
 sky130_fd_sc_hd__buf_2 _11544_ (.A(_06025_),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_4 _11545_ (.A(\CPU_Dmem_value_a5[15][17] ),
    .B(_06053_),
    .Y(_06063_));
 sky130_fd_sc_hd__a211o_4 _11546_ (.A1(_04721_),
    .A2(_06062_),
    .B1(_06050_),
    .C1(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__inv_2 _11547_ (.A(_06064_),
    .Y(_01055_));
 sky130_fd_sc_hd__buf_2 _11548_ (.A(_04660_),
    .X(_06065_));
 sky130_fd_sc_hd__nor2_4 _11549_ (.A(\CPU_Dmem_value_a5[15][16] ),
    .B(_06053_),
    .Y(_06066_));
 sky130_fd_sc_hd__a211o_4 _11550_ (.A1(_04725_),
    .A2(_06062_),
    .B1(_06065_),
    .C1(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__inv_2 _11551_ (.A(_06067_),
    .Y(_01054_));
 sky130_fd_sc_hd__buf_2 _11552_ (.A(_06024_),
    .X(_06068_));
 sky130_fd_sc_hd__nor2_4 _11553_ (.A(\CPU_Dmem_value_a5[15][15] ),
    .B(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__a211o_4 _11554_ (.A1(_04729_),
    .A2(_06062_),
    .B1(_06065_),
    .C1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__inv_2 _11555_ (.A(_06070_),
    .Y(_01053_));
 sky130_fd_sc_hd__nor2_4 _11556_ (.A(\CPU_Dmem_value_a5[15][14] ),
    .B(_06068_),
    .Y(_06071_));
 sky130_fd_sc_hd__a211o_4 _11557_ (.A1(_04733_),
    .A2(_06062_),
    .B1(_06065_),
    .C1(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__inv_2 _11558_ (.A(_06072_),
    .Y(_01052_));
 sky130_fd_sc_hd__nor2_4 _11559_ (.A(\CPU_Dmem_value_a5[15][13] ),
    .B(_06068_),
    .Y(_06073_));
 sky130_fd_sc_hd__a211o_4 _11560_ (.A1(_04739_),
    .A2(_06062_),
    .B1(_06065_),
    .C1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__inv_2 _11561_ (.A(_06074_),
    .Y(_01051_));
 sky130_fd_sc_hd__nor2_4 _11562_ (.A(\CPU_Dmem_value_a5[15][12] ),
    .B(_06068_),
    .Y(_06075_));
 sky130_fd_sc_hd__a211o_4 _11563_ (.A1(_04743_),
    .A2(_06062_),
    .B1(_06065_),
    .C1(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__inv_2 _11564_ (.A(_06076_),
    .Y(_01050_));
 sky130_fd_sc_hd__buf_2 _11565_ (.A(_06025_),
    .X(_06077_));
 sky130_fd_sc_hd__nor2_4 _11566_ (.A(\CPU_Dmem_value_a5[15][11] ),
    .B(_06068_),
    .Y(_06078_));
 sky130_fd_sc_hd__a211o_4 _11567_ (.A1(_04748_),
    .A2(_06077_),
    .B1(_06065_),
    .C1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__inv_2 _11568_ (.A(_06079_),
    .Y(_01049_));
 sky130_fd_sc_hd__buf_2 _11569_ (.A(_04660_),
    .X(_06080_));
 sky130_fd_sc_hd__nor2_4 _11570_ (.A(\CPU_Dmem_value_a5[15][10] ),
    .B(_06068_),
    .Y(_06081_));
 sky130_fd_sc_hd__a211o_4 _11571_ (.A1(_04752_),
    .A2(_06077_),
    .B1(_06080_),
    .C1(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__inv_2 _11572_ (.A(_06082_),
    .Y(_01048_));
 sky130_fd_sc_hd__buf_2 _11573_ (.A(_06024_),
    .X(_06083_));
 sky130_fd_sc_hd__nor2_4 _11574_ (.A(\CPU_Dmem_value_a5[15][9] ),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__a211o_4 _11575_ (.A1(_04756_),
    .A2(_06077_),
    .B1(_06080_),
    .C1(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__inv_2 _11576_ (.A(_06085_),
    .Y(_01047_));
 sky130_fd_sc_hd__nor2_4 _11577_ (.A(\CPU_Dmem_value_a5[15][8] ),
    .B(_06083_),
    .Y(_06086_));
 sky130_fd_sc_hd__a211o_4 _11578_ (.A1(_04760_),
    .A2(_06077_),
    .B1(_06080_),
    .C1(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__inv_2 _11579_ (.A(_06087_),
    .Y(_01046_));
 sky130_fd_sc_hd__nor2_4 _11580_ (.A(\CPU_Dmem_value_a5[15][7] ),
    .B(_06083_),
    .Y(_06088_));
 sky130_fd_sc_hd__a211o_4 _11581_ (.A1(_04766_),
    .A2(_06077_),
    .B1(_06080_),
    .C1(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__inv_2 _11582_ (.A(_06089_),
    .Y(_01045_));
 sky130_fd_sc_hd__nor2_4 _11583_ (.A(\CPU_Dmem_value_a5[15][6] ),
    .B(_06083_),
    .Y(_06090_));
 sky130_fd_sc_hd__a211o_4 _11584_ (.A1(_04770_),
    .A2(_06077_),
    .B1(_06080_),
    .C1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__inv_2 _11585_ (.A(_06091_),
    .Y(_01044_));
 sky130_fd_sc_hd__nor2_4 _11586_ (.A(\CPU_Dmem_value_a5[15][5] ),
    .B(_06083_),
    .Y(_06092_));
 sky130_fd_sc_hd__a211o_4 _11587_ (.A1(_04775_),
    .A2(_06027_),
    .B1(_06080_),
    .C1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__inv_2 _11588_ (.A(_06093_),
    .Y(_01043_));
 sky130_fd_sc_hd__nor2_4 _11589_ (.A(\CPU_Dmem_value_a5[15][4] ),
    .B(_06083_),
    .Y(_06094_));
 sky130_fd_sc_hd__a211o_4 _11590_ (.A1(_04779_),
    .A2(_06027_),
    .B1(_04888_),
    .C1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__inv_2 _11591_ (.A(_06095_),
    .Y(_01042_));
 sky130_fd_sc_hd__and2_4 _11592_ (.A(\CPU_Dmem_value_a5[15][3] ),
    .B(_06023_),
    .X(_06096_));
 sky130_fd_sc_hd__a211o_4 _11593_ (.A1(\CPU_dmem_wr_data_a4[3] ),
    .A2(_06026_),
    .B1(_05935_),
    .C1(_06096_),
    .X(_01041_));
 sky130_fd_sc_hd__and2_4 _11594_ (.A(\CPU_Dmem_value_a5[15][2] ),
    .B(_06023_),
    .X(_06097_));
 sky130_fd_sc_hd__a211o_4 _11595_ (.A1(\CPU_dmem_wr_data_a4[2] ),
    .A2(_06026_),
    .B1(_05935_),
    .C1(_06097_),
    .X(_01040_));
 sky130_fd_sc_hd__and2_4 _11596_ (.A(\CPU_Dmem_value_a5[15][1] ),
    .B(_06023_),
    .X(_06098_));
 sky130_fd_sc_hd__a211o_4 _11597_ (.A1(\CPU_dmem_wr_data_a4[1] ),
    .A2(_06026_),
    .B1(_04662_),
    .C1(_06098_),
    .X(_01039_));
 sky130_fd_sc_hd__and2_4 _11598_ (.A(\CPU_Dmem_value_a5[15][0] ),
    .B(_06023_),
    .X(_06099_));
 sky130_fd_sc_hd__a211o_4 _11599_ (.A1(\CPU_dmem_wr_data_a4[0] ),
    .A2(_06026_),
    .B1(_04662_),
    .C1(_06099_),
    .X(_01038_));
 sky130_fd_sc_hd__buf_2 _11600_ (.A(CPU_reset_a3),
    .X(_06100_));
 sky130_fd_sc_hd__buf_2 _11601_ (.A(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__buf_2 _11602_ (.A(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__buf_2 _11603_ (.A(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__buf_2 _11604_ (.A(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__inv_2 _11605_ (.A(\CPU_Xreg_value_a4[0][31] ),
    .Y(_06105_));
 sky130_fd_sc_hd__nor2_4 _11606_ (.A(_06104_),
    .B(_06105_),
    .Y(_01037_));
 sky130_fd_sc_hd__inv_2 _11607_ (.A(\CPU_Xreg_value_a4[0][30] ),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_4 _11608_ (.A(_06104_),
    .B(_06106_),
    .Y(_01036_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(\CPU_Xreg_value_a4[0][29] ),
    .Y(_06107_));
 sky130_fd_sc_hd__nor2_4 _11610_ (.A(_06104_),
    .B(_06107_),
    .Y(_01035_));
 sky130_fd_sc_hd__inv_2 _11611_ (.A(\CPU_Xreg_value_a4[0][28] ),
    .Y(_06108_));
 sky130_fd_sc_hd__nor2_4 _11612_ (.A(_06104_),
    .B(_06108_),
    .Y(_01034_));
 sky130_fd_sc_hd__inv_2 _11613_ (.A(\CPU_Xreg_value_a4[0][27] ),
    .Y(_06109_));
 sky130_fd_sc_hd__nor2_4 _11614_ (.A(_06104_),
    .B(_06109_),
    .Y(_01033_));
 sky130_fd_sc_hd__inv_2 _11615_ (.A(\CPU_Xreg_value_a4[0][26] ),
    .Y(_06110_));
 sky130_fd_sc_hd__nor2_4 _11616_ (.A(_06104_),
    .B(_06110_),
    .Y(_01032_));
 sky130_fd_sc_hd__buf_2 _11617_ (.A(_06103_),
    .X(_06111_));
 sky130_fd_sc_hd__inv_2 _11618_ (.A(\CPU_Xreg_value_a4[0][25] ),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_4 _11619_ (.A(_06111_),
    .B(_06112_),
    .Y(_01031_));
 sky130_fd_sc_hd__inv_2 _11620_ (.A(\CPU_Xreg_value_a4[0][24] ),
    .Y(_06113_));
 sky130_fd_sc_hd__nor2_4 _11621_ (.A(_06111_),
    .B(_06113_),
    .Y(_01030_));
 sky130_fd_sc_hd__inv_2 _11622_ (.A(\CPU_Xreg_value_a4[0][23] ),
    .Y(_06114_));
 sky130_fd_sc_hd__nor2_4 _11623_ (.A(_06111_),
    .B(_06114_),
    .Y(_01029_));
 sky130_fd_sc_hd__inv_2 _11624_ (.A(\CPU_Xreg_value_a4[0][22] ),
    .Y(_06115_));
 sky130_fd_sc_hd__nor2_4 _11625_ (.A(_06111_),
    .B(_06115_),
    .Y(_01028_));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(\CPU_Xreg_value_a4[0][21] ),
    .Y(_06116_));
 sky130_fd_sc_hd__nor2_4 _11627_ (.A(_06111_),
    .B(_06116_),
    .Y(_01027_));
 sky130_fd_sc_hd__inv_2 _11628_ (.A(\CPU_Xreg_value_a4[0][20] ),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_4 _11629_ (.A(_06111_),
    .B(_06117_),
    .Y(_01026_));
 sky130_fd_sc_hd__buf_2 _11630_ (.A(_06101_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_2 _11631_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__inv_2 _11632_ (.A(\CPU_Xreg_value_a4[0][19] ),
    .Y(_06120_));
 sky130_fd_sc_hd__nor2_4 _11633_ (.A(_06119_),
    .B(_06120_),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _11634_ (.A(\CPU_Xreg_value_a4[0][18] ),
    .Y(_06121_));
 sky130_fd_sc_hd__nor2_4 _11635_ (.A(_06119_),
    .B(_06121_),
    .Y(_01024_));
 sky130_fd_sc_hd__inv_2 _11636_ (.A(\CPU_Xreg_value_a4[0][17] ),
    .Y(_06122_));
 sky130_fd_sc_hd__nor2_4 _11637_ (.A(_06119_),
    .B(_06122_),
    .Y(_01023_));
 sky130_fd_sc_hd__inv_2 _11638_ (.A(\CPU_Xreg_value_a4[0][16] ),
    .Y(_06123_));
 sky130_fd_sc_hd__nor2_4 _11639_ (.A(_06119_),
    .B(_06123_),
    .Y(_01022_));
 sky130_fd_sc_hd__inv_2 _11640_ (.A(\CPU_Xreg_value_a4[0][15] ),
    .Y(_06124_));
 sky130_fd_sc_hd__nor2_4 _11641_ (.A(_06119_),
    .B(_06124_),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _11642_ (.A(\CPU_Xreg_value_a4[0][14] ),
    .Y(_06125_));
 sky130_fd_sc_hd__nor2_4 _11643_ (.A(_06119_),
    .B(_06125_),
    .Y(_01020_));
 sky130_fd_sc_hd__buf_2 _11644_ (.A(_06118_),
    .X(_06126_));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(\CPU_Xreg_value_a4[0][13] ),
    .Y(_06127_));
 sky130_fd_sc_hd__nor2_4 _11646_ (.A(_06126_),
    .B(_06127_),
    .Y(_01019_));
 sky130_fd_sc_hd__inv_2 _11647_ (.A(\CPU_Xreg_value_a4[0][12] ),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_4 _11648_ (.A(_06126_),
    .B(_06128_),
    .Y(_01018_));
 sky130_fd_sc_hd__inv_2 _11649_ (.A(\CPU_Xreg_value_a4[0][11] ),
    .Y(_06129_));
 sky130_fd_sc_hd__nor2_4 _11650_ (.A(_06126_),
    .B(_06129_),
    .Y(_01017_));
 sky130_fd_sc_hd__inv_2 _11651_ (.A(\CPU_Xreg_value_a4[0][10] ),
    .Y(_06130_));
 sky130_fd_sc_hd__nor2_4 _11652_ (.A(_06126_),
    .B(_06130_),
    .Y(_01016_));
 sky130_fd_sc_hd__inv_2 _11653_ (.A(\CPU_Xreg_value_a4[0][9] ),
    .Y(_06131_));
 sky130_fd_sc_hd__nor2_4 _11654_ (.A(_06126_),
    .B(_06131_),
    .Y(_01015_));
 sky130_fd_sc_hd__inv_2 _11655_ (.A(\CPU_Xreg_value_a4[0][8] ),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_4 _11656_ (.A(_06126_),
    .B(_06132_),
    .Y(_01014_));
 sky130_fd_sc_hd__buf_2 _11657_ (.A(_06118_),
    .X(_06133_));
 sky130_fd_sc_hd__inv_2 _11658_ (.A(\CPU_Xreg_value_a4[0][7] ),
    .Y(_06134_));
 sky130_fd_sc_hd__nor2_4 _11659_ (.A(_06133_),
    .B(_06134_),
    .Y(_01013_));
 sky130_fd_sc_hd__inv_2 _11660_ (.A(\CPU_Xreg_value_a4[0][6] ),
    .Y(_06135_));
 sky130_fd_sc_hd__nor2_4 _11661_ (.A(_06133_),
    .B(_06135_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _11662_ (.A(\CPU_Xreg_value_a4[0][5] ),
    .Y(_06136_));
 sky130_fd_sc_hd__nor2_4 _11663_ (.A(_06133_),
    .B(_06136_),
    .Y(_01011_));
 sky130_fd_sc_hd__inv_2 _11664_ (.A(\CPU_Xreg_value_a4[0][4] ),
    .Y(_06137_));
 sky130_fd_sc_hd__nor2_4 _11665_ (.A(_06133_),
    .B(_06137_),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _11666_ (.A(\CPU_Xreg_value_a4[0][3] ),
    .Y(_06138_));
 sky130_fd_sc_hd__nor2_4 _11667_ (.A(_06133_),
    .B(_06138_),
    .Y(_01009_));
 sky130_fd_sc_hd__inv_2 _11668_ (.A(\CPU_Xreg_value_a4[0][2] ),
    .Y(_06139_));
 sky130_fd_sc_hd__nor2_4 _11669_ (.A(_06133_),
    .B(_06139_),
    .Y(_01008_));
 sky130_fd_sc_hd__buf_2 _11670_ (.A(_06102_),
    .X(_06140_));
 sky130_fd_sc_hd__inv_2 _11671_ (.A(\CPU_Xreg_value_a4[0][1] ),
    .Y(_06141_));
 sky130_fd_sc_hd__nor2_4 _11672_ (.A(_06140_),
    .B(_06141_),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _11673_ (.A(\CPU_Xreg_value_a4[0][0] ),
    .Y(_06142_));
 sky130_fd_sc_hd__nor2_4 _11674_ (.A(_06140_),
    .B(_06142_),
    .Y(_01006_));
 sky130_fd_sc_hd__or4_4 _11675_ (.A(CPU_valid_load_a5),
    .B(CPU_valid_taken_br_a5),
    .C(CPU_valid_taken_br_a4),
    .D(\gen_clkP_CPU_dmem_rd_en_a5.pwr_en ),
    .X(_06143_));
 sky130_fd_sc_hd__inv_2 _11676_ (.A(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__o22a_4 _11677_ (.A1(\CPU_rd_a3[2] ),
    .A2(_06143_),
    .B1(\CPU_rd_a5[2] ),
    .B2(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__buf_2 _11678_ (.A(_06143_),
    .X(_06146_));
 sky130_fd_sc_hd__o22a_4 _11679_ (.A1(\CPU_rd_a3[3] ),
    .A2(_06146_),
    .B1(\CPU_rd_a5[3] ),
    .B2(_06144_),
    .X(_06147_));
 sky130_fd_sc_hd__or2_4 _11680_ (.A(_06145_),
    .B(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__o22a_4 _11681_ (.A1(\CPU_rd_a3[0] ),
    .A2(_06146_),
    .B1(\CPU_rd_a5[0] ),
    .B2(_06144_),
    .X(_06149_));
 sky130_fd_sc_hd__inv_2 _11682_ (.A(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__o22a_4 _11683_ (.A1(\CPU_rd_a3[1] ),
    .A2(_06146_),
    .B1(\CPU_rd_a5[1] ),
    .B2(_06144_),
    .X(_06151_));
 sky130_fd_sc_hd__or2_4 _11684_ (.A(_06150_),
    .B(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__or2_4 _11685_ (.A(_06148_),
    .B(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__buf_2 _11686_ (.A(_06144_),
    .X(_06154_));
 sky130_fd_sc_hd__o22a_4 _11687_ (.A1(\CPU_rd_a3[4] ),
    .A2(_06146_),
    .B1(\CPU_rd_a5[4] ),
    .B2(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__or2_4 _11688_ (.A(_06149_),
    .B(_06151_),
    .X(_06156_));
 sky130_fd_sc_hd__or2_4 _11689_ (.A(_06148_),
    .B(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__or2_4 _11690_ (.A(\CPU_rd_a3[0] ),
    .B(\CPU_rd_a3[1] ),
    .X(_06158_));
 sky130_fd_sc_hd__or4_4 _11691_ (.A(\CPU_rd_a3[2] ),
    .B(\CPU_rd_a3[3] ),
    .C(\CPU_rd_a3[4] ),
    .D(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__and3_4 _11692_ (.A(\gen_clkP_CPU_rd_valid_a4.pwr_en ),
    .B(_06144_),
    .C(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__or2_4 _11693_ (.A(CPU_valid_load_a5),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__buf_2 _11694_ (.A(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__o21ai_4 _11695_ (.A1(_06155_),
    .A2(_06157_),
    .B1(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__or2_4 _11696_ (.A(_06155_),
    .B(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__buf_2 _11697_ (.A(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__buf_2 _11698_ (.A(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__nor2_4 _11699_ (.A(_06153_),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__buf_2 _11700_ (.A(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__buf_2 _11701_ (.A(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__buf_2 _11702_ (.A(_06154_),
    .X(_06170_));
 sky130_fd_sc_hd__buf_2 _11703_ (.A(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__buf_2 _11704_ (.A(_06146_),
    .X(_06172_));
 sky130_fd_sc_hd__buf_2 _11705_ (.A(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__inv_2 _11706_ (.A(CPU_is_addi_a3),
    .Y(_06174_));
 sky130_fd_sc_hd__or3_4 _11707_ (.A(CPU_is_slti_a3),
    .B(CPU_is_slt_a3),
    .C(CPU_is_add_a3),
    .X(_06175_));
 sky130_fd_sc_hd__and2_4 _11708_ (.A(_06174_),
    .B(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__buf_2 _11709_ (.A(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__inv_2 _11710_ (.A(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__buf_2 _11711_ (.A(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__buf_2 _11712_ (.A(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__inv_2 _11713_ (.A(\CPU_src1_value_a3[30] ),
    .Y(_06181_));
 sky130_fd_sc_hd__inv_2 _11714_ (.A(\CPU_imm_a3[10] ),
    .Y(_06182_));
 sky130_fd_sc_hd__buf_2 _11715_ (.A(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__buf_2 _11716_ (.A(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__buf_2 _11717_ (.A(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__buf_2 _11718_ (.A(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__buf_2 _11719_ (.A(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__buf_2 _11720_ (.A(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__buf_2 _11721_ (.A(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__buf_2 _11722_ (.A(\CPU_imm_a3[10] ),
    .X(_06190_));
 sky130_fd_sc_hd__buf_2 _11723_ (.A(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__buf_2 _11724_ (.A(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__buf_2 _11725_ (.A(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__buf_2 _11726_ (.A(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__buf_2 _11727_ (.A(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__o22a_4 _11728_ (.A1(_06181_),
    .A2(_06188_),
    .B1(\CPU_src1_value_a3[30] ),
    .B2(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__inv_2 _11729_ (.A(\CPU_src1_value_a3[29] ),
    .Y(_06197_));
 sky130_fd_sc_hd__o22a_4 _11730_ (.A1(_06197_),
    .A2(_06186_),
    .B1(\CPU_src1_value_a3[29] ),
    .B2(_06194_),
    .X(_06198_));
 sky130_fd_sc_hd__inv_2 _11731_ (.A(\CPU_src1_value_a3[28] ),
    .Y(_06199_));
 sky130_fd_sc_hd__buf_2 _11732_ (.A(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__o22a_4 _11733_ (.A1(_06200_),
    .A2(_06188_),
    .B1(\CPU_src1_value_a3[28] ),
    .B2(_06195_),
    .X(_06201_));
 sky130_fd_sc_hd__and2_4 _11734_ (.A(\CPU_src1_value_a3[27] ),
    .B(_06193_),
    .X(_06202_));
 sky130_fd_sc_hd__and2_4 _11735_ (.A(\CPU_src1_value_a3[26] ),
    .B(_06193_),
    .X(_06203_));
 sky130_fd_sc_hd__inv_2 _11736_ (.A(\CPU_src1_value_a3[25] ),
    .Y(_06204_));
 sky130_fd_sc_hd__inv_2 _11737_ (.A(\CPU_src1_value_a3[24] ),
    .Y(_06205_));
 sky130_fd_sc_hd__buf_2 _11738_ (.A(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__o22a_4 _11739_ (.A1(_06204_),
    .A2(_06188_),
    .B1(_06206_),
    .B2(_06188_),
    .X(_06207_));
 sky130_fd_sc_hd__inv_2 _11740_ (.A(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__inv_2 _11741_ (.A(\CPU_src1_value_a3[27] ),
    .Y(_06209_));
 sky130_fd_sc_hd__a21o_4 _11742_ (.A1(_06209_),
    .A2(_06186_),
    .B1(_06202_),
    .X(_06210_));
 sky130_fd_sc_hd__inv_2 _11743_ (.A(\CPU_src1_value_a3[26] ),
    .Y(_06211_));
 sky130_fd_sc_hd__a21o_4 _11744_ (.A1(_06211_),
    .A2(_06187_),
    .B1(_06203_),
    .X(_06212_));
 sky130_fd_sc_hd__o22a_4 _11745_ (.A1(_06204_),
    .A2(_06186_),
    .B1(\CPU_src1_value_a3[25] ),
    .B2(_06194_),
    .X(_06213_));
 sky130_fd_sc_hd__o22a_4 _11746_ (.A1(_06206_),
    .A2(_06187_),
    .B1(\CPU_src1_value_a3[24] ),
    .B2(_06194_),
    .X(_06214_));
 sky130_fd_sc_hd__nand2_4 _11747_ (.A(_06213_),
    .B(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__inv_2 _11748_ (.A(\CPU_src1_value_a3[21] ),
    .Y(_06216_));
 sky130_fd_sc_hd__inv_2 _11749_ (.A(\CPU_src1_value_a3[20] ),
    .Y(_06217_));
 sky130_fd_sc_hd__buf_2 _11750_ (.A(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__o22a_4 _11751_ (.A1(_06216_),
    .A2(_06186_),
    .B1(_06218_),
    .B2(_06186_),
    .X(_06219_));
 sky130_fd_sc_hd__inv_2 _11752_ (.A(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__inv_2 _11753_ (.A(\CPU_src1_value_a3[23] ),
    .Y(_06221_));
 sky130_fd_sc_hd__a2bb2o_4 _11754_ (.A1_N(_06221_),
    .A2_N(_06187_),
    .B1(\CPU_src1_value_a3[22] ),
    .B2(_06194_),
    .X(_06222_));
 sky130_fd_sc_hd__and2_4 _11755_ (.A(\CPU_src1_value_a3[17] ),
    .B(_06192_),
    .X(_06223_));
 sky130_fd_sc_hd__and2_4 _11756_ (.A(\CPU_src1_value_a3[16] ),
    .B(_06191_),
    .X(_06224_));
 sky130_fd_sc_hd__and2_4 _11757_ (.A(\CPU_src1_value_a3[19] ),
    .B(_06192_),
    .X(_06225_));
 sky130_fd_sc_hd__and2_4 _11758_ (.A(\CPU_src1_value_a3[18] ),
    .B(_06192_),
    .X(_06226_));
 sky130_fd_sc_hd__or4_4 _11759_ (.A(_06223_),
    .B(_06224_),
    .C(_06225_),
    .D(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__inv_2 _11760_ (.A(\CPU_src1_value_a3[13] ),
    .Y(_06228_));
 sky130_fd_sc_hd__buf_2 _11761_ (.A(_06184_),
    .X(_06229_));
 sky130_fd_sc_hd__inv_2 _11762_ (.A(\CPU_src1_value_a3[12] ),
    .Y(_06230_));
 sky130_fd_sc_hd__o22a_4 _11763_ (.A1(_06228_),
    .A2(_06229_),
    .B1(_06230_),
    .B2(_06229_),
    .X(_06231_));
 sky130_fd_sc_hd__inv_2 _11764_ (.A(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__inv_2 _11765_ (.A(\CPU_src1_value_a3[15] ),
    .Y(_06233_));
 sky130_fd_sc_hd__a2bb2o_4 _11766_ (.A1_N(_06233_),
    .A2_N(_06185_),
    .B1(\CPU_src1_value_a3[14] ),
    .B2(_06192_),
    .X(_06234_));
 sky130_fd_sc_hd__o22a_4 _11767_ (.A1(_06228_),
    .A2(_06184_),
    .B1(\CPU_src1_value_a3[13] ),
    .B2(_06190_),
    .X(_06235_));
 sky130_fd_sc_hd__inv_2 _11768_ (.A(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__o22a_4 _11769_ (.A1(_06230_),
    .A2(_06183_),
    .B1(\CPU_src1_value_a3[12] ),
    .B2(_06190_),
    .X(_06237_));
 sky130_fd_sc_hd__inv_2 _11770_ (.A(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__o22a_4 _11771_ (.A1(_06233_),
    .A2(_06183_),
    .B1(\CPU_src1_value_a3[15] ),
    .B2(_06190_),
    .X(_06239_));
 sky130_fd_sc_hd__inv_2 _11772_ (.A(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__inv_2 _11773_ (.A(\CPU_src1_value_a3[14] ),
    .Y(_06241_));
 sky130_fd_sc_hd__o22a_4 _11774_ (.A1(_06241_),
    .A2(_06184_),
    .B1(\CPU_src1_value_a3[14] ),
    .B2(_06190_),
    .X(_06242_));
 sky130_fd_sc_hd__inv_2 _11775_ (.A(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__or4_4 _11776_ (.A(_06236_),
    .B(_06238_),
    .C(_06240_),
    .D(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__or2_4 _11777_ (.A(\CPU_src1_value_a3[11] ),
    .B(\CPU_imm_a3[11] ),
    .X(_06245_));
 sky130_fd_sc_hd__and3_4 _11778_ (.A(\CPU_src1_value_a3[10] ),
    .B(_06191_),
    .C(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__a21bo_4 _11779_ (.A1(\CPU_src1_value_a3[11] ),
    .A2(\CPU_imm_a3[11] ),
    .B1_N(_06245_),
    .X(_06247_));
 sky130_fd_sc_hd__inv_2 _11780_ (.A(\CPU_src1_value_a3[10] ),
    .Y(_06248_));
 sky130_fd_sc_hd__o22a_4 _11781_ (.A1(_06248_),
    .A2(_06183_),
    .B1(\CPU_src1_value_a3[10] ),
    .B2(_06190_),
    .X(_06249_));
 sky130_fd_sc_hd__inv_2 _11782_ (.A(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__inv_2 _11783_ (.A(\CPU_src1_value_a3[9] ),
    .Y(_06251_));
 sky130_fd_sc_hd__inv_2 _11784_ (.A(\CPU_src1_value_a3[8] ),
    .Y(_06252_));
 sky130_fd_sc_hd__buf_2 _11785_ (.A(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__o22a_4 _11786_ (.A1(_06251_),
    .A2(_06183_),
    .B1(_06253_),
    .B2(_06183_),
    .X(_06254_));
 sky130_fd_sc_hd__or3_4 _11787_ (.A(_06247_),
    .B(_06250_),
    .C(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__inv_2 _11788_ (.A(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__a211o_4 _11789_ (.A1(\CPU_src1_value_a3[11] ),
    .A2(\CPU_imm_a3[11] ),
    .B1(_06246_),
    .C1(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__inv_2 _11790_ (.A(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__nor2_4 _11791_ (.A(_06244_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__o22a_4 _11792_ (.A1(_06251_),
    .A2(_06184_),
    .B1(\CPU_src1_value_a3[9] ),
    .B2(_06191_),
    .X(_06260_));
 sky130_fd_sc_hd__inv_2 _11793_ (.A(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__o22a_4 _11794_ (.A1(_06253_),
    .A2(_06184_),
    .B1(\CPU_src1_value_a3[8] ),
    .B2(_06191_),
    .X(_06262_));
 sky130_fd_sc_hd__inv_2 _11795_ (.A(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__or4_4 _11796_ (.A(_06247_),
    .B(_06250_),
    .C(_06261_),
    .D(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__inv_2 _11797_ (.A(\CPU_src1_value_a3[3] ),
    .Y(_06265_));
 sky130_fd_sc_hd__inv_2 _11798_ (.A(\CPU_imm_a3[3] ),
    .Y(_06266_));
 sky130_fd_sc_hd__inv_2 _11799_ (.A(\CPU_src1_value_a3[2] ),
    .Y(_06267_));
 sky130_fd_sc_hd__inv_2 _11800_ (.A(\CPU_imm_a3[2] ),
    .Y(_06268_));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(\CPU_src1_value_a3[1] ),
    .Y(_06269_));
 sky130_fd_sc_hd__inv_2 _11802_ (.A(\CPU_imm_a3[1] ),
    .Y(_06270_));
 sky130_fd_sc_hd__inv_2 _11803_ (.A(\CPU_src1_value_a3[0] ),
    .Y(_06271_));
 sky130_fd_sc_hd__inv_2 _11804_ (.A(\CPU_imm_a3[0] ),
    .Y(_06272_));
 sky130_fd_sc_hd__o22a_4 _11805_ (.A1(\CPU_src1_value_a3[1] ),
    .A2(_06270_),
    .B1(_06269_),
    .B2(\CPU_imm_a3[1] ),
    .X(_06273_));
 sky130_fd_sc_hd__or3_4 _11806_ (.A(_06271_),
    .B(_06272_),
    .C(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__o21a_4 _11807_ (.A1(_06269_),
    .A2(_06270_),
    .B1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__o22a_4 _11808_ (.A1(\CPU_src1_value_a3[2] ),
    .A2(_06268_),
    .B1(_06267_),
    .B2(\CPU_imm_a3[2] ),
    .X(_06276_));
 sky130_fd_sc_hd__or2_4 _11809_ (.A(_06275_),
    .B(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__o21a_4 _11810_ (.A1(_06267_),
    .A2(_06268_),
    .B1(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__o22a_4 _11811_ (.A1(\CPU_src1_value_a3[3] ),
    .A2(_06266_),
    .B1(_06265_),
    .B2(\CPU_imm_a3[3] ),
    .X(_06279_));
 sky130_fd_sc_hd__or2_4 _11812_ (.A(_06278_),
    .B(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__o21a_4 _11813_ (.A1(_06265_),
    .A2(_06266_),
    .B1(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__inv_2 _11814_ (.A(\CPU_src1_value_a3[7] ),
    .Y(_06282_));
 sky130_fd_sc_hd__o22a_4 _11815_ (.A1(_06282_),
    .A2(_06182_),
    .B1(\CPU_src1_value_a3[7] ),
    .B2(\CPU_imm_a3[10] ),
    .X(_06283_));
 sky130_fd_sc_hd__inv_2 _11816_ (.A(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__inv_2 _11817_ (.A(\CPU_src1_value_a3[6] ),
    .Y(_06285_));
 sky130_fd_sc_hd__o22a_4 _11818_ (.A1(_06285_),
    .A2(_06182_),
    .B1(\CPU_src1_value_a3[6] ),
    .B2(\CPU_imm_a3[10] ),
    .X(_06286_));
 sky130_fd_sc_hd__inv_2 _11819_ (.A(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__inv_2 _11820_ (.A(\CPU_src1_value_a3[5] ),
    .Y(_06288_));
 sky130_fd_sc_hd__or2_4 _11821_ (.A(_06288_),
    .B(_06182_),
    .X(_06289_));
 sky130_fd_sc_hd__inv_2 _11822_ (.A(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__or2_4 _11823_ (.A(\CPU_src1_value_a3[5] ),
    .B(\CPU_imm_a3[10] ),
    .X(_06291_));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__or2_4 _11825_ (.A(_06290_),
    .B(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__inv_2 _11826_ (.A(\CPU_src1_value_a3[4] ),
    .Y(_06294_));
 sky130_fd_sc_hd__and2_4 _11827_ (.A(_06294_),
    .B(\CPU_imm_a3[4] ),
    .X(_06295_));
 sky130_fd_sc_hd__or2_4 _11828_ (.A(_06294_),
    .B(\CPU_imm_a3[4] ),
    .X(_06296_));
 sky130_fd_sc_hd__inv_2 _11829_ (.A(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nor2_4 _11830_ (.A(_06295_),
    .B(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__or4_4 _11831_ (.A(_06284_),
    .B(_06287_),
    .C(_06293_),
    .D(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__or2_4 _11832_ (.A(\CPU_src1_value_a3[7] ),
    .B(\CPU_src1_value_a3[6] ),
    .X(_06300_));
 sky130_fd_sc_hd__and2_4 _11833_ (.A(\CPU_src1_value_a3[4] ),
    .B(\CPU_imm_a3[4] ),
    .X(_06301_));
 sky130_fd_sc_hd__or2_4 _11834_ (.A(_06290_),
    .B(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__and4_4 _11835_ (.A(_06283_),
    .B(_06286_),
    .C(_06291_),
    .D(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__a21oi_4 _11836_ (.A1(_06191_),
    .A2(_06300_),
    .B1(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__o21a_4 _11837_ (.A1(_06281_),
    .A2(_06299_),
    .B1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__or3_4 _11838_ (.A(_06264_),
    .B(_06244_),
    .C(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__inv_2 _11839_ (.A(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__or4_4 _11840_ (.A(_06232_),
    .B(_06234_),
    .C(_06259_),
    .D(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__inv_2 _11841_ (.A(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__o22a_4 _11842_ (.A1(_06221_),
    .A2(_06185_),
    .B1(\CPU_src1_value_a3[23] ),
    .B2(_06192_),
    .X(_06310_));
 sky130_fd_sc_hd__inv_2 _11843_ (.A(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__inv_2 _11844_ (.A(\CPU_src1_value_a3[22] ),
    .Y(_06312_));
 sky130_fd_sc_hd__o22a_4 _11845_ (.A1(_06312_),
    .A2(_06185_),
    .B1(\CPU_src1_value_a3[22] ),
    .B2(_06193_),
    .X(_06313_));
 sky130_fd_sc_hd__inv_2 _11846_ (.A(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__o22a_4 _11847_ (.A1(_06216_),
    .A2(_06185_),
    .B1(\CPU_src1_value_a3[21] ),
    .B2(_06193_),
    .X(_06315_));
 sky130_fd_sc_hd__o22a_4 _11848_ (.A1(_06217_),
    .A2(_06185_),
    .B1(\CPU_src1_value_a3[20] ),
    .B2(_06193_),
    .X(_06316_));
 sky130_fd_sc_hd__nand2_4 _11849_ (.A(_06315_),
    .B(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(\CPU_src1_value_a3[17] ),
    .Y(_06318_));
 sky130_fd_sc_hd__a21o_4 _11851_ (.A1(_06318_),
    .A2(_06229_),
    .B1(_06223_),
    .X(_06319_));
 sky130_fd_sc_hd__inv_2 _11852_ (.A(\CPU_src1_value_a3[16] ),
    .Y(_06320_));
 sky130_fd_sc_hd__a21o_4 _11853_ (.A1(_06320_),
    .A2(_06229_),
    .B1(_06224_),
    .X(_06321_));
 sky130_fd_sc_hd__inv_2 _11854_ (.A(\CPU_src1_value_a3[19] ),
    .Y(_06322_));
 sky130_fd_sc_hd__a21o_4 _11855_ (.A1(_06322_),
    .A2(_06229_),
    .B1(_06225_),
    .X(_06323_));
 sky130_fd_sc_hd__inv_2 _11856_ (.A(\CPU_src1_value_a3[18] ),
    .Y(_06324_));
 sky130_fd_sc_hd__a21o_4 _11857_ (.A1(_06324_),
    .A2(_06229_),
    .B1(_06226_),
    .X(_06325_));
 sky130_fd_sc_hd__or4_4 _11858_ (.A(_06319_),
    .B(_06321_),
    .C(_06323_),
    .D(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__or4_4 _11859_ (.A(_06311_),
    .B(_06314_),
    .C(_06317_),
    .D(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_4 _11860_ (.A(_06309_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__or4_4 _11861_ (.A(_06220_),
    .B(_06222_),
    .C(_06227_),
    .D(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__inv_2 _11862_ (.A(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__or4_4 _11863_ (.A(_06210_),
    .B(_06212_),
    .C(_06215_),
    .D(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__inv_2 _11864_ (.A(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__or4_4 _11865_ (.A(_06202_),
    .B(_06203_),
    .C(_06208_),
    .D(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__or2_4 _11866_ (.A(\CPU_src1_value_a3[29] ),
    .B(\CPU_src1_value_a3[28] ),
    .X(_06334_));
 sky130_fd_sc_hd__a32o_4 _11867_ (.A1(_06198_),
    .A2(_06201_),
    .A3(_06333_),
    .B1(_06195_),
    .B2(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__nand2_4 _11868_ (.A(_06196_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__o21a_4 _11869_ (.A1(_06181_),
    .A2(_06189_),
    .B1(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__inv_2 _11870_ (.A(\CPU_src1_value_a3[31] ),
    .Y(_06338_));
 sky130_fd_sc_hd__and2_4 _11871_ (.A(\CPU_src1_value_a3[31] ),
    .B(_06187_),
    .X(_06339_));
 sky130_fd_sc_hd__a21o_4 _11872_ (.A1(_06338_),
    .A2(_06195_),
    .B1(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__inv_2 _11873_ (.A(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__or2_4 _11874_ (.A(_06337_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nand2_4 _11875_ (.A(_06337_),
    .B(_06341_),
    .Y(_06343_));
 sky130_fd_sc_hd__inv_2 _11876_ (.A(\CPU_src2_value_a3[30] ),
    .Y(_06344_));
 sky130_fd_sc_hd__and2_4 _11877_ (.A(\CPU_src2_value_a3[30] ),
    .B(_06181_),
    .X(_06345_));
 sky130_fd_sc_hd__a21oi_4 _11878_ (.A1(_06344_),
    .A2(\CPU_src1_value_a3[30] ),
    .B1(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_4 _11879_ (.A(\CPU_src2_value_a3[29] ),
    .B(\CPU_src1_value_a3[29] ),
    .Y(_06347_));
 sky130_fd_sc_hd__inv_2 _11880_ (.A(\CPU_src2_value_a3[28] ),
    .Y(_06348_));
 sky130_fd_sc_hd__or2_4 _11881_ (.A(\CPU_src2_value_a3[29] ),
    .B(\CPU_src1_value_a3[29] ),
    .X(_06349_));
 sky130_fd_sc_hd__inv_2 _11882_ (.A(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__or3_4 _11883_ (.A(_06200_),
    .B(_06348_),
    .C(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__and2_4 _11884_ (.A(_06347_),
    .B(_06349_),
    .X(_06352_));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__o22a_4 _11886_ (.A1(_06200_),
    .A2(\CPU_src2_value_a3[28] ),
    .B1(\CPU_src1_value_a3[28] ),
    .B2(_06348_),
    .X(_06354_));
 sky130_fd_sc_hd__inv_2 _11887_ (.A(\CPU_src2_value_a3[27] ),
    .Y(_06355_));
 sky130_fd_sc_hd__or2_4 _11888_ (.A(_06355_),
    .B(_06209_),
    .X(_06356_));
 sky130_fd_sc_hd__inv_2 _11889_ (.A(\CPU_src2_value_a3[26] ),
    .Y(_06357_));
 sky130_fd_sc_hd__or2_4 _11890_ (.A(\CPU_src2_value_a3[27] ),
    .B(\CPU_src1_value_a3[27] ),
    .X(_06358_));
 sky130_fd_sc_hd__inv_2 _11891_ (.A(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__or3_4 _11892_ (.A(_06357_),
    .B(_06211_),
    .C(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__inv_2 _11893_ (.A(\CPU_src2_value_a3[25] ),
    .Y(_06361_));
 sky130_fd_sc_hd__or2_4 _11894_ (.A(_06361_),
    .B(_06204_),
    .X(_06362_));
 sky130_fd_sc_hd__inv_2 _11895_ (.A(\CPU_src2_value_a3[24] ),
    .Y(_06363_));
 sky130_fd_sc_hd__or2_4 _11896_ (.A(_06206_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__and2_4 _11897_ (.A(_06361_),
    .B(_06204_),
    .X(_06365_));
 sky130_fd_sc_hd__and2_4 _11898_ (.A(_06356_),
    .B(_06358_),
    .X(_06366_));
 sky130_fd_sc_hd__inv_2 _11899_ (.A(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__and2_4 _11900_ (.A(\CPU_src2_value_a3[26] ),
    .B(_06211_),
    .X(_06368_));
 sky130_fd_sc_hd__a21oi_4 _11901_ (.A1(_06357_),
    .A2(\CPU_src1_value_a3[26] ),
    .B1(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__or2_4 _11902_ (.A(_06367_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__a211o_4 _11903_ (.A1(_06362_),
    .A2(_06364_),
    .B1(_06365_),
    .C1(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__inv_2 _11904_ (.A(_06362_),
    .Y(_06372_));
 sky130_fd_sc_hd__or2_4 _11905_ (.A(_06372_),
    .B(_06365_),
    .X(_06373_));
 sky130_fd_sc_hd__o22a_4 _11906_ (.A1(_06206_),
    .A2(\CPU_src2_value_a3[24] ),
    .B1(\CPU_src1_value_a3[24] ),
    .B2(_06363_),
    .X(_06374_));
 sky130_fd_sc_hd__or2_4 _11907_ (.A(\CPU_src2_value_a3[23] ),
    .B(\CPU_src1_value_a3[23] ),
    .X(_06375_));
 sky130_fd_sc_hd__a21bo_4 _11908_ (.A1(\CPU_src2_value_a3[23] ),
    .A2(\CPU_src1_value_a3[23] ),
    .B1_N(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__inv_2 _11909_ (.A(\CPU_src2_value_a3[22] ),
    .Y(_06377_));
 sky130_fd_sc_hd__and2_4 _11910_ (.A(\CPU_src2_value_a3[22] ),
    .B(_06312_),
    .X(_06378_));
 sky130_fd_sc_hd__a21oi_4 _11911_ (.A1(_06377_),
    .A2(\CPU_src1_value_a3[22] ),
    .B1(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__inv_2 _11912_ (.A(\CPU_src2_value_a3[21] ),
    .Y(_06380_));
 sky130_fd_sc_hd__and2_4 _11913_ (.A(_06380_),
    .B(_06216_),
    .X(_06381_));
 sky130_fd_sc_hd__inv_2 _11914_ (.A(\CPU_src2_value_a3[20] ),
    .Y(_06382_));
 sky130_fd_sc_hd__o22a_4 _11915_ (.A1(_06380_),
    .A2(_06216_),
    .B1(_06218_),
    .B2(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__or4_4 _11916_ (.A(_06376_),
    .B(_06379_),
    .C(_06381_),
    .D(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__a32o_4 _11917_ (.A1(\CPU_src2_value_a3[22] ),
    .A2(\CPU_src1_value_a3[22] ),
    .A3(_06375_),
    .B1(\CPU_src2_value_a3[23] ),
    .B2(\CPU_src1_value_a3[23] ),
    .X(_06385_));
 sky130_fd_sc_hd__inv_2 _11918_ (.A(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__o22a_4 _11919_ (.A1(_06217_),
    .A2(\CPU_src2_value_a3[20] ),
    .B1(\CPU_src1_value_a3[20] ),
    .B2(_06382_),
    .X(_06387_));
 sky130_fd_sc_hd__a21o_4 _11920_ (.A1(\CPU_src2_value_a3[21] ),
    .A2(\CPU_src1_value_a3[21] ),
    .B1(_06381_),
    .X(_06388_));
 sky130_fd_sc_hd__or4_4 _11921_ (.A(_06376_),
    .B(_06379_),
    .C(_06387_),
    .D(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__inv_2 _11922_ (.A(\CPU_src2_value_a3[19] ),
    .Y(_06390_));
 sky130_fd_sc_hd__or2_4 _11923_ (.A(_06390_),
    .B(_06322_),
    .X(_06391_));
 sky130_fd_sc_hd__inv_2 _11924_ (.A(\CPU_src2_value_a3[18] ),
    .Y(_06392_));
 sky130_fd_sc_hd__or2_4 _11925_ (.A(\CPU_src2_value_a3[19] ),
    .B(\CPU_src1_value_a3[19] ),
    .X(_06393_));
 sky130_fd_sc_hd__inv_2 _11926_ (.A(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__or3_4 _11927_ (.A(_06392_),
    .B(_06324_),
    .C(_06394_),
    .X(_06395_));
 sky130_fd_sc_hd__nand2_4 _11928_ (.A(_06391_),
    .B(_06393_),
    .Y(_06396_));
 sky130_fd_sc_hd__or2_4 _11929_ (.A(_06392_),
    .B(\CPU_src1_value_a3[18] ),
    .X(_06397_));
 sky130_fd_sc_hd__o21a_4 _11930_ (.A1(\CPU_src2_value_a3[18] ),
    .A2(_06324_),
    .B1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__inv_2 _11931_ (.A(\CPU_src2_value_a3[17] ),
    .Y(_06399_));
 sky130_fd_sc_hd__and2_4 _11932_ (.A(_06399_),
    .B(_06318_),
    .X(_06400_));
 sky130_fd_sc_hd__inv_2 _11933_ (.A(\CPU_src2_value_a3[16] ),
    .Y(_06401_));
 sky130_fd_sc_hd__o22a_4 _11934_ (.A1(_06399_),
    .A2(_06318_),
    .B1(_06320_),
    .B2(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__or4_4 _11935_ (.A(_06396_),
    .B(_06398_),
    .C(_06400_),
    .D(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__and3_4 _11936_ (.A(_06391_),
    .B(_06395_),
    .C(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__or2_4 _11937_ (.A(_06389_),
    .B(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__o22a_4 _11938_ (.A1(_06320_),
    .A2(\CPU_src2_value_a3[16] ),
    .B1(\CPU_src1_value_a3[16] ),
    .B2(_06401_),
    .X(_06406_));
 sky130_fd_sc_hd__a21o_4 _11939_ (.A1(\CPU_src2_value_a3[17] ),
    .A2(\CPU_src1_value_a3[17] ),
    .B1(_06400_),
    .X(_06407_));
 sky130_fd_sc_hd__or4_4 _11940_ (.A(_06396_),
    .B(_06398_),
    .C(_06406_),
    .D(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__or2_4 _11941_ (.A(\CPU_src2_value_a3[15] ),
    .B(\CPU_src1_value_a3[15] ),
    .X(_06409_));
 sky130_fd_sc_hd__a21bo_4 _11942_ (.A1(\CPU_src2_value_a3[15] ),
    .A2(\CPU_src1_value_a3[15] ),
    .B1_N(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__inv_2 _11943_ (.A(\CPU_src2_value_a3[14] ),
    .Y(_06411_));
 sky130_fd_sc_hd__and2_4 _11944_ (.A(_06411_),
    .B(\CPU_src1_value_a3[14] ),
    .X(_06412_));
 sky130_fd_sc_hd__and2_4 _11945_ (.A(\CPU_src2_value_a3[14] ),
    .B(_06241_),
    .X(_06413_));
 sky130_fd_sc_hd__nor2_4 _11946_ (.A(_06412_),
    .B(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(\CPU_src2_value_a3[13] ),
    .Y(_06415_));
 sky130_fd_sc_hd__and2_4 _11948_ (.A(_06415_),
    .B(_06228_),
    .X(_06416_));
 sky130_fd_sc_hd__inv_2 _11949_ (.A(\CPU_src2_value_a3[12] ),
    .Y(_06417_));
 sky130_fd_sc_hd__o22a_4 _11950_ (.A1(_06415_),
    .A2(_06228_),
    .B1(_06230_),
    .B2(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__or4_4 _11951_ (.A(_06410_),
    .B(_06414_),
    .C(_06416_),
    .D(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__a32o_4 _11952_ (.A1(\CPU_src2_value_a3[14] ),
    .A2(\CPU_src1_value_a3[14] ),
    .A3(_06409_),
    .B1(\CPU_src2_value_a3[15] ),
    .B2(\CPU_src1_value_a3[15] ),
    .X(_06420_));
 sky130_fd_sc_hd__inv_2 _11953_ (.A(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__o22a_4 _11954_ (.A1(_06230_),
    .A2(\CPU_src2_value_a3[12] ),
    .B1(\CPU_src1_value_a3[12] ),
    .B2(_06417_),
    .X(_06422_));
 sky130_fd_sc_hd__a21o_4 _11955_ (.A1(\CPU_src2_value_a3[13] ),
    .A2(\CPU_src1_value_a3[13] ),
    .B1(_06416_),
    .X(_06423_));
 sky130_fd_sc_hd__or4_4 _11956_ (.A(_06410_),
    .B(_06414_),
    .C(_06422_),
    .D(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__nand2_4 _11957_ (.A(\CPU_src2_value_a3[11] ),
    .B(\CPU_src1_value_a3[11] ),
    .Y(_06425_));
 sky130_fd_sc_hd__inv_2 _11958_ (.A(\CPU_src2_value_a3[10] ),
    .Y(_06426_));
 sky130_fd_sc_hd__or2_4 _11959_ (.A(\CPU_src2_value_a3[11] ),
    .B(\CPU_src1_value_a3[11] ),
    .X(_06427_));
 sky130_fd_sc_hd__inv_2 _11960_ (.A(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__or3_4 _11961_ (.A(_06426_),
    .B(_06248_),
    .C(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__and2_4 _11962_ (.A(_06425_),
    .B(_06427_),
    .X(_06430_));
 sky130_fd_sc_hd__inv_2 _11963_ (.A(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__and2_4 _11964_ (.A(_06426_),
    .B(\CPU_src1_value_a3[10] ),
    .X(_06432_));
 sky130_fd_sc_hd__and2_4 _11965_ (.A(\CPU_src2_value_a3[10] ),
    .B(_06248_),
    .X(_06433_));
 sky130_fd_sc_hd__nor2_4 _11966_ (.A(_06432_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__inv_2 _11967_ (.A(\CPU_src2_value_a3[9] ),
    .Y(_06435_));
 sky130_fd_sc_hd__and2_4 _11968_ (.A(_06435_),
    .B(_06251_),
    .X(_06436_));
 sky130_fd_sc_hd__inv_2 _11969_ (.A(\CPU_src2_value_a3[8] ),
    .Y(_06437_));
 sky130_fd_sc_hd__o22a_4 _11970_ (.A1(_06435_),
    .A2(_06251_),
    .B1(_06252_),
    .B2(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__or4_4 _11971_ (.A(_06431_),
    .B(_06434_),
    .C(_06436_),
    .D(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__and3_4 _11972_ (.A(_06425_),
    .B(_06429_),
    .C(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__or2_4 _11973_ (.A(_06424_),
    .B(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__o22a_4 _11974_ (.A1(_06253_),
    .A2(\CPU_src2_value_a3[8] ),
    .B1(\CPU_src1_value_a3[8] ),
    .B2(_06437_),
    .X(_06442_));
 sky130_fd_sc_hd__a21o_4 _11975_ (.A1(\CPU_src2_value_a3[9] ),
    .A2(\CPU_src1_value_a3[9] ),
    .B1(_06436_),
    .X(_06443_));
 sky130_fd_sc_hd__or4_4 _11976_ (.A(_06431_),
    .B(_06434_),
    .C(_06442_),
    .D(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__nand2_4 _11977_ (.A(\CPU_src2_value_a3[7] ),
    .B(\CPU_src1_value_a3[7] ),
    .Y(_06445_));
 sky130_fd_sc_hd__inv_2 _11978_ (.A(\CPU_src2_value_a3[6] ),
    .Y(_06446_));
 sky130_fd_sc_hd__or2_4 _11979_ (.A(\CPU_src2_value_a3[7] ),
    .B(\CPU_src1_value_a3[7] ),
    .X(_06447_));
 sky130_fd_sc_hd__inv_2 _11980_ (.A(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__or3_4 _11981_ (.A(_06446_),
    .B(_06285_),
    .C(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__inv_2 _11982_ (.A(\CPU_src2_value_a3[5] ),
    .Y(_06450_));
 sky130_fd_sc_hd__or2_4 _11983_ (.A(_06450_),
    .B(_06288_),
    .X(_06451_));
 sky130_fd_sc_hd__inv_2 _11984_ (.A(\CPU_src2_value_a3[4] ),
    .Y(_06452_));
 sky130_fd_sc_hd__or2_4 _11985_ (.A(_06294_),
    .B(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__and2_4 _11986_ (.A(_06450_),
    .B(_06288_),
    .X(_06454_));
 sky130_fd_sc_hd__and2_4 _11987_ (.A(_06445_),
    .B(_06447_),
    .X(_06455_));
 sky130_fd_sc_hd__inv_2 _11988_ (.A(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__and2_4 _11989_ (.A(\CPU_src2_value_a3[6] ),
    .B(_06285_),
    .X(_06457_));
 sky130_fd_sc_hd__a21oi_4 _11990_ (.A1(_06446_),
    .A2(\CPU_src1_value_a3[6] ),
    .B1(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__or2_4 _11991_ (.A(_06456_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__a211o_4 _11992_ (.A1(_06451_),
    .A2(_06453_),
    .B1(_06454_),
    .C1(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__inv_2 _11993_ (.A(_06451_),
    .Y(_06461_));
 sky130_fd_sc_hd__or2_4 _11994_ (.A(_06461_),
    .B(_06454_),
    .X(_06462_));
 sky130_fd_sc_hd__o22a_4 _11995_ (.A1(_06294_),
    .A2(\CPU_src2_value_a3[4] ),
    .B1(\CPU_src1_value_a3[4] ),
    .B2(_06452_),
    .X(_06463_));
 sky130_fd_sc_hd__inv_2 _11996_ (.A(\CPU_src2_value_a3[3] ),
    .Y(_06464_));
 sky130_fd_sc_hd__and2_4 _11997_ (.A(_06464_),
    .B(_06265_),
    .X(_06465_));
 sky130_fd_sc_hd__inv_2 _11998_ (.A(\CPU_src2_value_a3[2] ),
    .Y(_06466_));
 sky130_fd_sc_hd__and2_4 _11999_ (.A(_06466_),
    .B(_06267_),
    .X(_06467_));
 sky130_fd_sc_hd__inv_2 _12000_ (.A(\CPU_src2_value_a3[1] ),
    .Y(_06468_));
 sky130_fd_sc_hd__inv_2 _12001_ (.A(\CPU_src2_value_a3[0] ),
    .Y(_06469_));
 sky130_fd_sc_hd__or2_4 _12002_ (.A(_06469_),
    .B(_06271_),
    .X(_06470_));
 sky130_fd_sc_hd__or2_4 _12003_ (.A(_06468_),
    .B(\CPU_src1_value_a3[1] ),
    .X(_06471_));
 sky130_fd_sc_hd__o21a_4 _12004_ (.A1(\CPU_src2_value_a3[1] ),
    .A2(_06269_),
    .B1(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__or2_4 _12005_ (.A(_06470_),
    .B(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__o21a_4 _12006_ (.A1(_06468_),
    .A2(_06269_),
    .B1(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__o22a_4 _12007_ (.A1(_06466_),
    .A2(_06267_),
    .B1(_06467_),
    .B2(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__o22a_4 _12008_ (.A1(_06464_),
    .A2(_06265_),
    .B1(_06465_),
    .B2(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__or4_4 _12009_ (.A(_06462_),
    .B(_06463_),
    .C(_06459_),
    .D(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__and4_4 _12010_ (.A(_06445_),
    .B(_06449_),
    .C(_06460_),
    .D(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__or3_4 _12011_ (.A(_06424_),
    .B(_06444_),
    .C(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__and4_4 _12012_ (.A(_06419_),
    .B(_06421_),
    .C(_06441_),
    .D(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__or3_4 _12013_ (.A(_06408_),
    .B(_06389_),
    .C(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__and4_4 _12014_ (.A(_06384_),
    .B(_06386_),
    .C(_06405_),
    .D(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__or4_4 _12015_ (.A(_06373_),
    .B(_06374_),
    .C(_06370_),
    .D(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__and4_4 _12016_ (.A(_06356_),
    .B(_06360_),
    .C(_06371_),
    .D(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__or3_4 _12017_ (.A(_06353_),
    .B(_06354_),
    .C(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__and3_4 _12018_ (.A(_06347_),
    .B(_06351_),
    .C(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__or2_4 _12019_ (.A(_06346_),
    .B(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__o21a_4 _12020_ (.A1(_06344_),
    .A2(_06181_),
    .B1(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__or2_4 _12021_ (.A(_06338_),
    .B(\CPU_src2_value_a3[31] ),
    .X(_06489_));
 sky130_fd_sc_hd__inv_2 _12022_ (.A(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__and2_4 _12023_ (.A(_06338_),
    .B(\CPU_src2_value_a3[31] ),
    .X(_06491_));
 sky130_fd_sc_hd__or2_4 _12024_ (.A(_06490_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__inv_2 _12025_ (.A(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_4 _12026_ (.A(_06488_),
    .B(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__inv_2 _12027_ (.A(CPU_is_add_a3),
    .Y(_06495_));
 sky130_fd_sc_hd__or2_4 _12028_ (.A(_06495_),
    .B(CPU_is_addi_a3),
    .X(_06496_));
 sky130_fd_sc_hd__buf_2 _12029_ (.A(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__inv_2 _12030_ (.A(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__buf_2 _12031_ (.A(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__o21a_4 _12032_ (.A1(_06488_),
    .A2(_06493_),
    .B1(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__a32o_4 _12033_ (.A1(_06180_),
    .A2(_06342_),
    .A3(_06343_),
    .B1(_06494_),
    .B2(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__o22a_4 _12034_ (.A1(\CPU_dmem_rd_data_a5[31] ),
    .A2(_06171_),
    .B1(_06173_),
    .B2(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__inv_2 _12035_ (.A(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__buf_2 _12036_ (.A(_06168_),
    .X(_06504_));
 sky130_fd_sc_hd__nor2_4 _12037_ (.A(\CPU_Xreg_value_a4[1][31] ),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__a211o_4 _12038_ (.A1(_06169_),
    .A2(_06503_),
    .B1(_06118_),
    .C1(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__inv_2 _12039_ (.A(_06506_),
    .Y(_01005_));
 sky130_fd_sc_hd__buf_2 _12040_ (.A(_06172_),
    .X(_06507_));
 sky130_fd_sc_hd__buf_2 _12041_ (.A(_06498_),
    .X(_06508_));
 sky130_fd_sc_hd__buf_2 _12042_ (.A(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2_4 _12043_ (.A(_06346_),
    .B(_06486_),
    .Y(_06510_));
 sky130_fd_sc_hd__or2_4 _12044_ (.A(_06196_),
    .B(_06335_),
    .X(_06511_));
 sky130_fd_sc_hd__and2_4 _12045_ (.A(_06336_),
    .B(_06178_),
    .X(_06512_));
 sky130_fd_sc_hd__a32o_4 _12046_ (.A1(_06487_),
    .A2(_06509_),
    .A3(_06510_),
    .B1(_06511_),
    .B2(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__o22a_4 _12047_ (.A1(\CPU_dmem_rd_data_a5[30] ),
    .A2(_06171_),
    .B1(_06507_),
    .B2(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__inv_2 _12048_ (.A(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__nor2_4 _12049_ (.A(\CPU_Xreg_value_a4[1][30] ),
    .B(_06504_),
    .Y(_06516_));
 sky130_fd_sc_hd__a211o_4 _12050_ (.A1(_06169_),
    .A2(_06515_),
    .B1(_06118_),
    .C1(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__inv_2 _12051_ (.A(_06517_),
    .Y(_01004_));
 sky130_fd_sc_hd__inv_2 _12052_ (.A(_06198_),
    .Y(_06518_));
 sky130_fd_sc_hd__buf_2 _12053_ (.A(_06189_),
    .X(_06519_));
 sky130_fd_sc_hd__nand2_4 _12054_ (.A(_06333_),
    .B(_06201_),
    .Y(_06520_));
 sky130_fd_sc_hd__o21a_4 _12055_ (.A1(_06200_),
    .A2(_06519_),
    .B1(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__or2_4 _12056_ (.A(_06518_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__nand2_4 _12057_ (.A(_06518_),
    .B(_06521_),
    .Y(_06523_));
 sky130_fd_sc_hd__or2_4 _12058_ (.A(_06484_),
    .B(_06354_),
    .X(_06524_));
 sky130_fd_sc_hd__o21a_4 _12059_ (.A1(_06200_),
    .A2(_06348_),
    .B1(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__or2_4 _12060_ (.A(_06353_),
    .B(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__buf_2 _12061_ (.A(_06497_),
    .X(_06527_));
 sky130_fd_sc_hd__a21oi_4 _12062_ (.A1(_06353_),
    .A2(_06525_),
    .B1(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__a32o_4 _12063_ (.A1(_06180_),
    .A2(_06522_),
    .A3(_06523_),
    .B1(_06526_),
    .B2(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__o22a_4 _12064_ (.A1(\CPU_dmem_rd_data_a5[29] ),
    .A2(_06171_),
    .B1(_06507_),
    .B2(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__inv_2 _12065_ (.A(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__nor2_4 _12066_ (.A(\CPU_Xreg_value_a4[1][29] ),
    .B(_06504_),
    .Y(_06532_));
 sky130_fd_sc_hd__a211o_4 _12067_ (.A1(_06169_),
    .A2(_06531_),
    .B1(_06118_),
    .C1(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__inv_2 _12068_ (.A(_06533_),
    .Y(_01003_));
 sky130_fd_sc_hd__or2_4 _12069_ (.A(_06333_),
    .B(_06201_),
    .X(_06534_));
 sky130_fd_sc_hd__nand2_4 _12070_ (.A(_06484_),
    .B(_06354_),
    .Y(_06535_));
 sky130_fd_sc_hd__and2_4 _12071_ (.A(_06508_),
    .B(_06524_),
    .X(_06536_));
 sky130_fd_sc_hd__a32o_4 _12072_ (.A1(_06180_),
    .A2(_06520_),
    .A3(_06534_),
    .B1(_06535_),
    .B2(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__o22a_4 _12073_ (.A1(\CPU_dmem_rd_data_a5[28] ),
    .A2(_06171_),
    .B1(_06507_),
    .B2(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__inv_2 _12074_ (.A(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__buf_2 _12075_ (.A(_06102_),
    .X(_06540_));
 sky130_fd_sc_hd__buf_2 _12076_ (.A(_06168_),
    .X(_06541_));
 sky130_fd_sc_hd__nor2_4 _12077_ (.A(\CPU_Xreg_value_a4[1][28] ),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__a211o_4 _12078_ (.A1(_06169_),
    .A2(_06539_),
    .B1(_06540_),
    .C1(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__inv_2 _12079_ (.A(_06543_),
    .Y(_01002_));
 sky130_fd_sc_hd__buf_2 _12080_ (.A(_06167_),
    .X(_06544_));
 sky130_fd_sc_hd__buf_2 _12081_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_2 _12082_ (.A(_06179_),
    .X(_06546_));
 sky130_fd_sc_hd__inv_2 _12083_ (.A(_06210_),
    .Y(_06547_));
 sky130_fd_sc_hd__o21a_4 _12084_ (.A1(_06330_),
    .A2(_06215_),
    .B1(_06207_),
    .X(_06548_));
 sky130_fd_sc_hd__nor2_4 _12085_ (.A(_06212_),
    .B(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__or2_4 _12086_ (.A(_06203_),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__nand2_4 _12087_ (.A(_06547_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__or2_4 _12088_ (.A(_06547_),
    .B(_06550_),
    .X(_06552_));
 sky130_fd_sc_hd__inv_2 _12089_ (.A(_06364_),
    .Y(_06553_));
 sky130_fd_sc_hd__nor2_4 _12090_ (.A(_06482_),
    .B(_06374_),
    .Y(_06554_));
 sky130_fd_sc_hd__or2_4 _12091_ (.A(_06553_),
    .B(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__inv_2 _12092_ (.A(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__o21a_4 _12093_ (.A1(_06365_),
    .A2(_06556_),
    .B1(_06362_),
    .X(_06557_));
 sky130_fd_sc_hd__or2_4 _12094_ (.A(_06369_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__o21a_4 _12095_ (.A1(_06357_),
    .A2(_06211_),
    .B1(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__or2_4 _12096_ (.A(_06367_),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__a21oi_4 _12097_ (.A1(_06367_),
    .A2(_06559_),
    .B1(_06527_),
    .Y(_06561_));
 sky130_fd_sc_hd__a32o_4 _12098_ (.A1(_06546_),
    .A2(_06551_),
    .A3(_06552_),
    .B1(_06560_),
    .B2(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__o22a_4 _12099_ (.A1(\CPU_dmem_rd_data_a5[27] ),
    .A2(_06171_),
    .B1(_06507_),
    .B2(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__inv_2 _12100_ (.A(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__nor2_4 _12101_ (.A(\CPU_Xreg_value_a4[1][27] ),
    .B(_06541_),
    .Y(_06565_));
 sky130_fd_sc_hd__a211o_4 _12102_ (.A1(_06545_),
    .A2(_06564_),
    .B1(_06540_),
    .C1(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__inv_2 _12103_ (.A(_06566_),
    .Y(_01001_));
 sky130_fd_sc_hd__buf_2 _12104_ (.A(_06154_),
    .X(_06567_));
 sky130_fd_sc_hd__a211o_4 _12105_ (.A1(_06212_),
    .A2(_06548_),
    .B1(_06177_),
    .C1(_06549_),
    .X(_06568_));
 sky130_fd_sc_hd__inv_2 _12106_ (.A(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__nand2_4 _12107_ (.A(_06369_),
    .B(_06557_),
    .Y(_06570_));
 sky130_fd_sc_hd__and3_4 _12108_ (.A(_06499_),
    .B(_06558_),
    .C(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__or2_4 _12109_ (.A(_06569_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__o22a_4 _12110_ (.A1(\CPU_dmem_rd_data_a5[26] ),
    .A2(_06567_),
    .B1(_06507_),
    .B2(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__inv_2 _12111_ (.A(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__nor2_4 _12112_ (.A(\CPU_Xreg_value_a4[1][26] ),
    .B(_06541_),
    .Y(_06575_));
 sky130_fd_sc_hd__a211o_4 _12113_ (.A1(_06545_),
    .A2(_06574_),
    .B1(_06540_),
    .C1(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__inv_2 _12114_ (.A(_06576_),
    .Y(_01000_));
 sky130_fd_sc_hd__buf_2 _12115_ (.A(_06499_),
    .X(_06577_));
 sky130_fd_sc_hd__or2_4 _12116_ (.A(_06373_),
    .B(_06556_),
    .X(_06578_));
 sky130_fd_sc_hd__inv_2 _12117_ (.A(_06373_),
    .Y(_06579_));
 sky130_fd_sc_hd__or2_4 _12118_ (.A(_06579_),
    .B(_06555_),
    .X(_06580_));
 sky130_fd_sc_hd__buf_2 _12119_ (.A(_06178_),
    .X(_06581_));
 sky130_fd_sc_hd__buf_2 _12120_ (.A(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__inv_2 _12121_ (.A(_06214_),
    .Y(_06583_));
 sky130_fd_sc_hd__or2_4 _12122_ (.A(_06330_),
    .B(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__o21a_4 _12123_ (.A1(_06206_),
    .A2(_06519_),
    .B1(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__a2bb2o_4 _12124_ (.A1_N(_06213_),
    .A2_N(_06585_),
    .B1(_06213_),
    .B2(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__a32o_4 _12125_ (.A1(_06577_),
    .A2(_06578_),
    .A3(_06580_),
    .B1(_06582_),
    .B2(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__o22a_4 _12126_ (.A1(\CPU_dmem_rd_data_a5[25] ),
    .A2(_06567_),
    .B1(_06507_),
    .B2(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__inv_2 _12127_ (.A(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__nor2_4 _12128_ (.A(\CPU_Xreg_value_a4[1][25] ),
    .B(_06541_),
    .Y(_06590_));
 sky130_fd_sc_hd__a211o_4 _12129_ (.A1(_06545_),
    .A2(_06589_),
    .B1(_06540_),
    .C1(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__inv_2 _12130_ (.A(_06591_),
    .Y(_00999_));
 sky130_fd_sc_hd__buf_2 _12131_ (.A(_06172_),
    .X(_06592_));
 sky130_fd_sc_hd__or2_4 _12132_ (.A(_06329_),
    .B(_06214_),
    .X(_06593_));
 sky130_fd_sc_hd__and3_4 _12133_ (.A(_06179_),
    .B(_06584_),
    .C(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__a211o_4 _12134_ (.A1(_06482_),
    .A2(_06374_),
    .B1(_06497_),
    .C1(_06554_),
    .X(_06595_));
 sky130_fd_sc_hd__inv_2 _12135_ (.A(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__or2_4 _12136_ (.A(_06594_),
    .B(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__o22a_4 _12137_ (.A1(\CPU_dmem_rd_data_a5[24] ),
    .A2(_06567_),
    .B1(_06592_),
    .B2(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__inv_2 _12138_ (.A(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__nor2_4 _12139_ (.A(\CPU_Xreg_value_a4[1][24] ),
    .B(_06541_),
    .Y(_06600_));
 sky130_fd_sc_hd__a211o_4 _12140_ (.A1(_06545_),
    .A2(_06599_),
    .B1(_06540_),
    .C1(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__inv_2 _12141_ (.A(_06601_),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _12142_ (.A(_06227_),
    .Y(_06602_));
 sky130_fd_sc_hd__o21a_4 _12143_ (.A1(_06309_),
    .A2(_06326_),
    .B1(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__o21a_4 _12144_ (.A1(_06317_),
    .A2(_06603_),
    .B1(_06219_),
    .X(_06604_));
 sky130_fd_sc_hd__or2_4 _12145_ (.A(_06314_),
    .B(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__o21a_4 _12146_ (.A1(_06312_),
    .A2(_06519_),
    .B1(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__or2_4 _12147_ (.A(_06311_),
    .B(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_4 _12148_ (.A(_06311_),
    .B(_06606_),
    .Y(_06608_));
 sky130_fd_sc_hd__o21a_4 _12149_ (.A1(_06480_),
    .A2(_06408_),
    .B1(_06404_),
    .X(_06609_));
 sky130_fd_sc_hd__or2_4 _12150_ (.A(_06387_),
    .B(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__o21a_4 _12151_ (.A1(_06218_),
    .A2(_06382_),
    .B1(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__o22a_4 _12152_ (.A1(_06380_),
    .A2(_06216_),
    .B1(_06381_),
    .B2(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__or2_4 _12153_ (.A(_06379_),
    .B(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__o21a_4 _12154_ (.A1(_06377_),
    .A2(_06312_),
    .B1(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__or2_4 _12155_ (.A(_06376_),
    .B(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__a21oi_4 _12156_ (.A1(_06376_),
    .A2(_06614_),
    .B1(_06527_),
    .Y(_06616_));
 sky130_fd_sc_hd__a32o_4 _12157_ (.A1(_06546_),
    .A2(_06607_),
    .A3(_06608_),
    .B1(_06615_),
    .B2(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__o22a_4 _12158_ (.A1(\CPU_dmem_rd_data_a5[23] ),
    .A2(_06567_),
    .B1(_06592_),
    .B2(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__inv_2 _12159_ (.A(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nor2_4 _12160_ (.A(\CPU_Xreg_value_a4[1][23] ),
    .B(_06541_),
    .Y(_06620_));
 sky130_fd_sc_hd__a211o_4 _12161_ (.A1(_06545_),
    .A2(_06619_),
    .B1(_06540_),
    .C1(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__inv_2 _12162_ (.A(_06621_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_4 _12163_ (.A(_06379_),
    .B(_06612_),
    .Y(_06622_));
 sky130_fd_sc_hd__nand2_4 _12164_ (.A(_06314_),
    .B(_06604_),
    .Y(_06623_));
 sky130_fd_sc_hd__and2_4 _12165_ (.A(_06179_),
    .B(_06605_),
    .X(_06624_));
 sky130_fd_sc_hd__a32o_4 _12166_ (.A1(_06577_),
    .A2(_06613_),
    .A3(_06622_),
    .B1(_06623_),
    .B2(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__o22a_4 _12167_ (.A1(\CPU_dmem_rd_data_a5[22] ),
    .A2(_06567_),
    .B1(_06592_),
    .B2(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__inv_2 _12168_ (.A(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__buf_2 _12169_ (.A(_06101_),
    .X(_06628_));
 sky130_fd_sc_hd__buf_2 _12170_ (.A(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__buf_2 _12171_ (.A(_06168_),
    .X(_06630_));
 sky130_fd_sc_hd__nor2_4 _12172_ (.A(\CPU_Xreg_value_a4[1][22] ),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__a211o_4 _12173_ (.A1(_06545_),
    .A2(_06627_),
    .B1(_06629_),
    .C1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__inv_2 _12174_ (.A(_06632_),
    .Y(_00996_));
 sky130_fd_sc_hd__buf_2 _12175_ (.A(_06544_),
    .X(_06633_));
 sky130_fd_sc_hd__or2_4 _12176_ (.A(_06388_),
    .B(_06611_),
    .X(_06634_));
 sky130_fd_sc_hd__nand2_4 _12177_ (.A(_06388_),
    .B(_06611_),
    .Y(_06635_));
 sky130_fd_sc_hd__inv_2 _12178_ (.A(_06316_),
    .Y(_06636_));
 sky130_fd_sc_hd__or2_4 _12179_ (.A(_06636_),
    .B(_06603_),
    .X(_06637_));
 sky130_fd_sc_hd__o21a_4 _12180_ (.A1(_06218_),
    .A2(_06519_),
    .B1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__a2bb2o_4 _12181_ (.A1_N(_06315_),
    .A2_N(_06638_),
    .B1(_06315_),
    .B2(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__a32o_4 _12182_ (.A1(_06577_),
    .A2(_06634_),
    .A3(_06635_),
    .B1(_06582_),
    .B2(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__o22a_4 _12183_ (.A1(\CPU_dmem_rd_data_a5[21] ),
    .A2(_06567_),
    .B1(_06592_),
    .B2(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__inv_2 _12184_ (.A(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nor2_4 _12185_ (.A(\CPU_Xreg_value_a4[1][21] ),
    .B(_06630_),
    .Y(_06643_));
 sky130_fd_sc_hd__a211o_4 _12186_ (.A1(_06633_),
    .A2(_06642_),
    .B1(_06629_),
    .C1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__inv_2 _12187_ (.A(_06644_),
    .Y(_00995_));
 sky130_fd_sc_hd__buf_2 _12188_ (.A(_06154_),
    .X(_06645_));
 sky130_fd_sc_hd__nand2_4 _12189_ (.A(_06636_),
    .B(_06603_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2_4 _12190_ (.A(_06387_),
    .B(_06609_),
    .Y(_06647_));
 sky130_fd_sc_hd__and2_4 _12191_ (.A(_06508_),
    .B(_06610_),
    .X(_06648_));
 sky130_fd_sc_hd__a32o_4 _12192_ (.A1(_06546_),
    .A2(_06637_),
    .A3(_06646_),
    .B1(_06647_),
    .B2(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__o22a_4 _12193_ (.A1(\CPU_dmem_rd_data_a5[20] ),
    .A2(_06645_),
    .B1(_06592_),
    .B2(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__inv_2 _12194_ (.A(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__nor2_4 _12195_ (.A(\CPU_Xreg_value_a4[1][20] ),
    .B(_06630_),
    .Y(_06652_));
 sky130_fd_sc_hd__a211o_4 _12196_ (.A1(_06633_),
    .A2(_06651_),
    .B1(_06629_),
    .C1(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__inv_2 _12197_ (.A(_06653_),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _12198_ (.A(_06323_),
    .Y(_06654_));
 sky130_fd_sc_hd__inv_2 _12199_ (.A(_06325_),
    .Y(_06655_));
 sky130_fd_sc_hd__inv_2 _12200_ (.A(_06319_),
    .Y(_06656_));
 sky130_fd_sc_hd__inv_2 _12201_ (.A(_06321_),
    .Y(_06657_));
 sky130_fd_sc_hd__and3_4 _12202_ (.A(_06656_),
    .B(_06657_),
    .C(_06308_),
    .X(_06658_));
 sky130_fd_sc_hd__or3_4 _12203_ (.A(_06223_),
    .B(_06224_),
    .C(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__and2_4 _12204_ (.A(_06655_),
    .B(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__or2_4 _12205_ (.A(_06226_),
    .B(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__nand2_4 _12206_ (.A(_06654_),
    .B(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__or2_4 _12207_ (.A(_06654_),
    .B(_06661_),
    .X(_06663_));
 sky130_fd_sc_hd__or2_4 _12208_ (.A(_06480_),
    .B(_06406_),
    .X(_06664_));
 sky130_fd_sc_hd__o21a_4 _12209_ (.A1(_06320_),
    .A2(_06401_),
    .B1(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__o22a_4 _12210_ (.A1(_06399_),
    .A2(_06318_),
    .B1(_06400_),
    .B2(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__or2_4 _12211_ (.A(_06398_),
    .B(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__o21a_4 _12212_ (.A1(_06392_),
    .A2(_06324_),
    .B1(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__or2_4 _12213_ (.A(_06396_),
    .B(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__a21oi_4 _12214_ (.A1(_06396_),
    .A2(_06668_),
    .B1(_06527_),
    .Y(_06670_));
 sky130_fd_sc_hd__a32o_4 _12215_ (.A1(_06546_),
    .A2(_06662_),
    .A3(_06663_),
    .B1(_06669_),
    .B2(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__o22a_4 _12216_ (.A1(\CPU_dmem_rd_data_a5[19] ),
    .A2(_06645_),
    .B1(_06592_),
    .B2(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__inv_2 _12217_ (.A(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_4 _12218_ (.A(\CPU_Xreg_value_a4[1][19] ),
    .B(_06630_),
    .Y(_06674_));
 sky130_fd_sc_hd__a211o_4 _12219_ (.A1(_06633_),
    .A2(_06673_),
    .B1(_06629_),
    .C1(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_06675_),
    .Y(_00993_));
 sky130_fd_sc_hd__buf_2 _12221_ (.A(_06172_),
    .X(_06676_));
 sky130_fd_sc_hd__nand2_4 _12222_ (.A(_06398_),
    .B(_06666_),
    .Y(_06677_));
 sky130_fd_sc_hd__or2_4 _12223_ (.A(_06655_),
    .B(_06659_),
    .X(_06678_));
 sky130_fd_sc_hd__nor2_4 _12224_ (.A(_06177_),
    .B(_06660_),
    .Y(_06679_));
 sky130_fd_sc_hd__a32o_4 _12225_ (.A1(_06577_),
    .A2(_06667_),
    .A3(_06677_),
    .B1(_06678_),
    .B2(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__o22a_4 _12226_ (.A1(\CPU_dmem_rd_data_a5[18] ),
    .A2(_06645_),
    .B1(_06676_),
    .B2(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__inv_2 _12227_ (.A(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__nor2_4 _12228_ (.A(\CPU_Xreg_value_a4[1][18] ),
    .B(_06630_),
    .Y(_06683_));
 sky130_fd_sc_hd__a211o_4 _12229_ (.A1(_06633_),
    .A2(_06682_),
    .B1(_06629_),
    .C1(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__inv_2 _12230_ (.A(_06684_),
    .Y(_00992_));
 sky130_fd_sc_hd__or2_4 _12231_ (.A(_06407_),
    .B(_06665_),
    .X(_06685_));
 sky130_fd_sc_hd__nand2_4 _12232_ (.A(_06407_),
    .B(_06665_),
    .Y(_06686_));
 sky130_fd_sc_hd__and2_4 _12233_ (.A(_06308_),
    .B(_06657_),
    .X(_06687_));
 sky130_fd_sc_hd__nor2_4 _12234_ (.A(_06224_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__a2bb2o_4 _12235_ (.A1_N(_06656_),
    .A2_N(_06688_),
    .B1(_06656_),
    .B2(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__a32o_4 _12236_ (.A1(_06577_),
    .A2(_06685_),
    .A3(_06686_),
    .B1(_06582_),
    .B2(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__o22a_4 _12237_ (.A1(\CPU_dmem_rd_data_a5[17] ),
    .A2(_06645_),
    .B1(_06676_),
    .B2(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__inv_2 _12238_ (.A(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__nor2_4 _12239_ (.A(\CPU_Xreg_value_a4[1][17] ),
    .B(_06630_),
    .Y(_06693_));
 sky130_fd_sc_hd__a211o_4 _12240_ (.A1(_06633_),
    .A2(_06692_),
    .B1(_06629_),
    .C1(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__inv_2 _12241_ (.A(_06694_),
    .Y(_00991_));
 sky130_fd_sc_hd__a211o_4 _12242_ (.A1(_06309_),
    .A2(_06321_),
    .B1(_06177_),
    .C1(_06687_),
    .X(_06695_));
 sky130_fd_sc_hd__inv_2 _12243_ (.A(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_4 _12244_ (.A(_06480_),
    .B(_06406_),
    .Y(_06697_));
 sky130_fd_sc_hd__and3_4 _12245_ (.A(_06499_),
    .B(_06664_),
    .C(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__or2_4 _12246_ (.A(_06696_),
    .B(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__o22a_4 _12247_ (.A1(\CPU_dmem_rd_data_a5[16] ),
    .A2(_06645_),
    .B1(_06676_),
    .B2(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__inv_2 _12248_ (.A(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__buf_2 _12249_ (.A(_06628_),
    .X(_06702_));
 sky130_fd_sc_hd__buf_2 _12250_ (.A(_06167_),
    .X(_06703_));
 sky130_fd_sc_hd__nor2_4 _12251_ (.A(\CPU_Xreg_value_a4[1][16] ),
    .B(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__a211o_4 _12252_ (.A1(_06633_),
    .A2(_06701_),
    .B1(_06702_),
    .C1(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__inv_2 _12253_ (.A(_06705_),
    .Y(_00990_));
 sky130_fd_sc_hd__buf_2 _12254_ (.A(_06168_),
    .X(_06706_));
 sky130_fd_sc_hd__o21a_4 _12255_ (.A1(_06305_),
    .A2(_06264_),
    .B1(_06258_),
    .X(_06707_));
 sky130_fd_sc_hd__or3_4 _12256_ (.A(_06236_),
    .B(_06238_),
    .C(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__and2_4 _12257_ (.A(_06231_),
    .B(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__or2_4 _12258_ (.A(_06243_),
    .B(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__o21a_4 _12259_ (.A1(_06241_),
    .A2(_06189_),
    .B1(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__or2_4 _12260_ (.A(_06240_),
    .B(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__nand2_4 _12261_ (.A(_06240_),
    .B(_06711_),
    .Y(_06713_));
 sky130_fd_sc_hd__o21a_4 _12262_ (.A1(_06478_),
    .A2(_06444_),
    .B1(_06440_),
    .X(_06714_));
 sky130_fd_sc_hd__or2_4 _12263_ (.A(_06422_),
    .B(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__o21a_4 _12264_ (.A1(_06230_),
    .A2(_06417_),
    .B1(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__o22a_4 _12265_ (.A1(_06415_),
    .A2(_06228_),
    .B1(_06416_),
    .B2(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__or2_4 _12266_ (.A(_06414_),
    .B(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__o21a_4 _12267_ (.A1(_06411_),
    .A2(_06241_),
    .B1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__or2_4 _12268_ (.A(_06410_),
    .B(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__a21oi_4 _12269_ (.A1(_06410_),
    .A2(_06719_),
    .B1(_06527_),
    .Y(_06721_));
 sky130_fd_sc_hd__a32o_4 _12270_ (.A1(_06546_),
    .A2(_06712_),
    .A3(_06713_),
    .B1(_06720_),
    .B2(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__o22a_4 _12271_ (.A1(\CPU_dmem_rd_data_a5[15] ),
    .A2(_06645_),
    .B1(_06676_),
    .B2(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__inv_2 _12272_ (.A(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__nor2_4 _12273_ (.A(\CPU_Xreg_value_a4[1][15] ),
    .B(_06703_),
    .Y(_06725_));
 sky130_fd_sc_hd__a211o_4 _12274_ (.A1(_06706_),
    .A2(_06724_),
    .B1(_06702_),
    .C1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__inv_2 _12275_ (.A(_06726_),
    .Y(_00989_));
 sky130_fd_sc_hd__buf_2 _12276_ (.A(_06154_),
    .X(_06727_));
 sky130_fd_sc_hd__nand2_4 _12277_ (.A(_06414_),
    .B(_06717_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand2_4 _12278_ (.A(_06243_),
    .B(_06709_),
    .Y(_06729_));
 sky130_fd_sc_hd__and2_4 _12279_ (.A(_06179_),
    .B(_06710_),
    .X(_06730_));
 sky130_fd_sc_hd__a32o_4 _12280_ (.A1(_06509_),
    .A2(_06718_),
    .A3(_06728_),
    .B1(_06729_),
    .B2(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__o22a_4 _12281_ (.A1(\CPU_dmem_rd_data_a5[14] ),
    .A2(_06727_),
    .B1(_06676_),
    .B2(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__inv_2 _12282_ (.A(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__nor2_4 _12283_ (.A(\CPU_Xreg_value_a4[1][14] ),
    .B(_06703_),
    .Y(_06734_));
 sky130_fd_sc_hd__a211o_4 _12284_ (.A1(_06706_),
    .A2(_06733_),
    .B1(_06702_),
    .C1(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__inv_2 _12285_ (.A(_06735_),
    .Y(_00988_));
 sky130_fd_sc_hd__or2_4 _12286_ (.A(_06423_),
    .B(_06716_),
    .X(_06736_));
 sky130_fd_sc_hd__nand2_4 _12287_ (.A(_06423_),
    .B(_06716_),
    .Y(_06737_));
 sky130_fd_sc_hd__or2_4 _12288_ (.A(_06238_),
    .B(_06707_),
    .X(_06738_));
 sky130_fd_sc_hd__o21a_4 _12289_ (.A1(_06230_),
    .A2(_06519_),
    .B1(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__a2bb2o_4 _12290_ (.A1_N(_06235_),
    .A2_N(_06739_),
    .B1(_06235_),
    .B2(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__a32o_4 _12291_ (.A1(_06509_),
    .A2(_06736_),
    .A3(_06737_),
    .B1(_06582_),
    .B2(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__o22a_4 _12292_ (.A1(\CPU_dmem_rd_data_a5[13] ),
    .A2(_06727_),
    .B1(_06676_),
    .B2(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__inv_2 _12293_ (.A(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_4 _12294_ (.A(\CPU_Xreg_value_a4[1][13] ),
    .B(_06703_),
    .Y(_06744_));
 sky130_fd_sc_hd__a211o_4 _12295_ (.A1(_06706_),
    .A2(_06743_),
    .B1(_06702_),
    .C1(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__inv_2 _12296_ (.A(_06745_),
    .Y(_00987_));
 sky130_fd_sc_hd__buf_2 _12297_ (.A(_06146_),
    .X(_06746_));
 sky130_fd_sc_hd__nand2_4 _12298_ (.A(_06238_),
    .B(_06707_),
    .Y(_06747_));
 sky130_fd_sc_hd__nand2_4 _12299_ (.A(_06422_),
    .B(_06714_),
    .Y(_06748_));
 sky130_fd_sc_hd__and2_4 _12300_ (.A(_06508_),
    .B(_06715_),
    .X(_06749_));
 sky130_fd_sc_hd__a32o_4 _12301_ (.A1(_06546_),
    .A2(_06738_),
    .A3(_06747_),
    .B1(_06748_),
    .B2(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__o22a_4 _12302_ (.A1(\CPU_dmem_rd_data_a5[12] ),
    .A2(_06727_),
    .B1(_06746_),
    .B2(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__inv_2 _12303_ (.A(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__nor2_4 _12304_ (.A(\CPU_Xreg_value_a4[1][12] ),
    .B(_06703_),
    .Y(_06753_));
 sky130_fd_sc_hd__a211o_4 _12305_ (.A1(_06706_),
    .A2(_06752_),
    .B1(_06702_),
    .C1(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__inv_2 _12306_ (.A(_06754_),
    .Y(_00986_));
 sky130_fd_sc_hd__or3_4 _12307_ (.A(_06261_),
    .B(_06263_),
    .C(_06305_),
    .X(_06755_));
 sky130_fd_sc_hd__and2_4 _12308_ (.A(_06254_),
    .B(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__or2_4 _12309_ (.A(_06250_),
    .B(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__o21a_4 _12310_ (.A1(_06248_),
    .A2(_06189_),
    .B1(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__or2_4 _12311_ (.A(_06247_),
    .B(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__nand2_4 _12312_ (.A(_06247_),
    .B(_06758_),
    .Y(_06760_));
 sky130_fd_sc_hd__or2_4 _12313_ (.A(_06478_),
    .B(_06442_),
    .X(_06761_));
 sky130_fd_sc_hd__o21a_4 _12314_ (.A1(_06253_),
    .A2(_06437_),
    .B1(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__o22a_4 _12315_ (.A1(_06435_),
    .A2(_06251_),
    .B1(_06436_),
    .B2(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__or2_4 _12316_ (.A(_06434_),
    .B(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__o21a_4 _12317_ (.A1(_06426_),
    .A2(_06248_),
    .B1(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__or2_4 _12318_ (.A(_06431_),
    .B(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__a21oi_4 _12319_ (.A1(_06431_),
    .A2(_06765_),
    .B1(_06527_),
    .Y(_06767_));
 sky130_fd_sc_hd__a32o_4 _12320_ (.A1(_06581_),
    .A2(_06759_),
    .A3(_06760_),
    .B1(_06766_),
    .B2(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__o22a_4 _12321_ (.A1(\CPU_dmem_rd_data_a5[11] ),
    .A2(_06727_),
    .B1(_06746_),
    .B2(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__inv_2 _12322_ (.A(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__nor2_4 _12323_ (.A(\CPU_Xreg_value_a4[1][11] ),
    .B(_06703_),
    .Y(_06771_));
 sky130_fd_sc_hd__a211o_4 _12324_ (.A1(_06706_),
    .A2(_06770_),
    .B1(_06702_),
    .C1(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__inv_2 _12325_ (.A(_06772_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_4 _12326_ (.A(_06434_),
    .B(_06763_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand2_4 _12327_ (.A(_06250_),
    .B(_06756_),
    .Y(_06774_));
 sky130_fd_sc_hd__and2_4 _12328_ (.A(_06179_),
    .B(_06757_),
    .X(_06775_));
 sky130_fd_sc_hd__a32o_4 _12329_ (.A1(_06509_),
    .A2(_06764_),
    .A3(_06773_),
    .B1(_06774_),
    .B2(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__o22a_4 _12330_ (.A1(\CPU_dmem_rd_data_a5[10] ),
    .A2(_06727_),
    .B1(_06746_),
    .B2(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__inv_2 _12331_ (.A(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__buf_2 _12332_ (.A(_06628_),
    .X(_06779_));
 sky130_fd_sc_hd__buf_2 _12333_ (.A(_06167_),
    .X(_06780_));
 sky130_fd_sc_hd__nor2_4 _12334_ (.A(\CPU_Xreg_value_a4[1][10] ),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__a211o_4 _12335_ (.A1(_06706_),
    .A2(_06778_),
    .B1(_06779_),
    .C1(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__inv_2 _12336_ (.A(_06782_),
    .Y(_00984_));
 sky130_fd_sc_hd__buf_2 _12337_ (.A(_06168_),
    .X(_06783_));
 sky130_fd_sc_hd__or2_4 _12338_ (.A(_06443_),
    .B(_06762_),
    .X(_06784_));
 sky130_fd_sc_hd__nand2_4 _12339_ (.A(_06443_),
    .B(_06762_),
    .Y(_06785_));
 sky130_fd_sc_hd__or2_4 _12340_ (.A(_06305_),
    .B(_06263_),
    .X(_06786_));
 sky130_fd_sc_hd__o21a_4 _12341_ (.A1(_06253_),
    .A2(_06519_),
    .B1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__a2bb2o_4 _12342_ (.A1_N(_06260_),
    .A2_N(_06787_),
    .B1(_06260_),
    .B2(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__a32o_4 _12343_ (.A1(_06509_),
    .A2(_06784_),
    .A3(_06785_),
    .B1(_06582_),
    .B2(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__o22a_4 _12344_ (.A1(\CPU_dmem_rd_data_a5[9] ),
    .A2(_06727_),
    .B1(_06746_),
    .B2(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__inv_2 _12345_ (.A(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__nor2_4 _12346_ (.A(\CPU_Xreg_value_a4[1][9] ),
    .B(_06780_),
    .Y(_06792_));
 sky130_fd_sc_hd__a211o_4 _12347_ (.A1(_06783_),
    .A2(_06791_),
    .B1(_06779_),
    .C1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__inv_2 _12348_ (.A(_06793_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_4 _12349_ (.A(_06305_),
    .B(_06263_),
    .Y(_06794_));
 sky130_fd_sc_hd__nand2_4 _12350_ (.A(_06478_),
    .B(_06442_),
    .Y(_06795_));
 sky130_fd_sc_hd__and2_4 _12351_ (.A(_06508_),
    .B(_06761_),
    .X(_06796_));
 sky130_fd_sc_hd__a32o_4 _12352_ (.A1(_06581_),
    .A2(_06786_),
    .A3(_06794_),
    .B1(_06795_),
    .B2(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__o22a_4 _12353_ (.A1(\CPU_dmem_rd_data_a5[8] ),
    .A2(_06170_),
    .B1(_06746_),
    .B2(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__inv_2 _12354_ (.A(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__nor2_4 _12355_ (.A(\CPU_Xreg_value_a4[1][8] ),
    .B(_06780_),
    .Y(_06800_));
 sky130_fd_sc_hd__a211o_4 _12356_ (.A1(_06783_),
    .A2(_06799_),
    .B1(_06779_),
    .C1(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__inv_2 _12357_ (.A(_06801_),
    .Y(_00982_));
 sky130_fd_sc_hd__nor2_4 _12358_ (.A(_06281_),
    .B(_06298_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_4 _12359_ (.A(_06301_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__o21a_4 _12360_ (.A1(_06292_),
    .A2(_06803_),
    .B1(_06289_),
    .X(_06804_));
 sky130_fd_sc_hd__or2_4 _12361_ (.A(_06287_),
    .B(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__o21a_4 _12362_ (.A1(_06285_),
    .A2(_06189_),
    .B1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__or2_4 _12363_ (.A(_06284_),
    .B(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__nand2_4 _12364_ (.A(_06284_),
    .B(_06806_),
    .Y(_06808_));
 sky130_fd_sc_hd__inv_2 _12365_ (.A(_06453_),
    .Y(_06809_));
 sky130_fd_sc_hd__nor2_4 _12366_ (.A(_06476_),
    .B(_06463_),
    .Y(_06810_));
 sky130_fd_sc_hd__or2_4 _12367_ (.A(_06809_),
    .B(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__inv_2 _12368_ (.A(_06811_),
    .Y(_06812_));
 sky130_fd_sc_hd__o21a_4 _12369_ (.A1(_06454_),
    .A2(_06812_),
    .B1(_06451_),
    .X(_06813_));
 sky130_fd_sc_hd__or2_4 _12370_ (.A(_06458_),
    .B(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__o21a_4 _12371_ (.A1(_06446_),
    .A2(_06285_),
    .B1(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__or2_4 _12372_ (.A(_06456_),
    .B(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__a21oi_4 _12373_ (.A1(_06456_),
    .A2(_06815_),
    .B1(_06497_),
    .Y(_06817_));
 sky130_fd_sc_hd__a32o_4 _12374_ (.A1(_06581_),
    .A2(_06807_),
    .A3(_06808_),
    .B1(_06816_),
    .B2(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__o22a_4 _12375_ (.A1(\CPU_dmem_rd_data_a5[7] ),
    .A2(_06170_),
    .B1(_06746_),
    .B2(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__inv_2 _12376_ (.A(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__nor2_4 _12377_ (.A(\CPU_Xreg_value_a4[1][7] ),
    .B(_06780_),
    .Y(_06821_));
 sky130_fd_sc_hd__a211o_4 _12378_ (.A1(_06783_),
    .A2(_06820_),
    .B1(_06779_),
    .C1(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__inv_2 _12379_ (.A(_06822_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_4 _12380_ (.A(_06287_),
    .B(_06804_),
    .Y(_06823_));
 sky130_fd_sc_hd__nand2_4 _12381_ (.A(_06458_),
    .B(_06813_),
    .Y(_06824_));
 sky130_fd_sc_hd__and2_4 _12382_ (.A(_06508_),
    .B(_06814_),
    .X(_06825_));
 sky130_fd_sc_hd__a32o_4 _12383_ (.A1(_06581_),
    .A2(_06805_),
    .A3(_06823_),
    .B1(_06824_),
    .B2(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__o22a_4 _12384_ (.A1(\CPU_dmem_rd_data_a5[6] ),
    .A2(_06170_),
    .B1(_06172_),
    .B2(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__inv_2 _12385_ (.A(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__nor2_4 _12386_ (.A(\CPU_Xreg_value_a4[1][6] ),
    .B(_06780_),
    .Y(_06829_));
 sky130_fd_sc_hd__a211o_4 _12387_ (.A1(_06783_),
    .A2(_06828_),
    .B1(_06779_),
    .C1(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__inv_2 _12388_ (.A(_06830_),
    .Y(_00980_));
 sky130_fd_sc_hd__or2_4 _12389_ (.A(_06462_),
    .B(_06812_),
    .X(_06831_));
 sky130_fd_sc_hd__inv_2 _12390_ (.A(_06462_),
    .Y(_06832_));
 sky130_fd_sc_hd__or2_4 _12391_ (.A(_06832_),
    .B(_06811_),
    .X(_06833_));
 sky130_fd_sc_hd__inv_2 _12392_ (.A(_06293_),
    .Y(_06834_));
 sky130_fd_sc_hd__a2bb2o_4 _12393_ (.A1_N(_06834_),
    .A2_N(_06803_),
    .B1(_06834_),
    .B2(_06803_),
    .X(_06835_));
 sky130_fd_sc_hd__a32o_4 _12394_ (.A1(_06509_),
    .A2(_06831_),
    .A3(_06833_),
    .B1(_06180_),
    .B2(_06835_),
    .X(\CPU_result_a3[5] ));
 sky130_fd_sc_hd__o22a_4 _12395_ (.A1(\CPU_dmem_rd_data_a5[5] ),
    .A2(_06170_),
    .B1(_06172_),
    .B2(\CPU_result_a3[5] ),
    .X(_06836_));
 sky130_fd_sc_hd__inv_2 _12396_ (.A(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__nor2_4 _12397_ (.A(\CPU_Xreg_value_a4[1][5] ),
    .B(_06780_),
    .Y(_06838_));
 sky130_fd_sc_hd__a211o_4 _12398_ (.A1(_06783_),
    .A2(_06837_),
    .B1(_06779_),
    .C1(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__inv_2 _12399_ (.A(_06839_),
    .Y(_00979_));
 sky130_fd_sc_hd__buf_2 _12400_ (.A(_06170_),
    .X(CPU_valid_a3));
 sky130_fd_sc_hd__a211o_4 _12401_ (.A1(_06281_),
    .A2(_06298_),
    .B1(_06177_),
    .C1(_06802_),
    .X(_06840_));
 sky130_fd_sc_hd__a211o_4 _12402_ (.A1(_06476_),
    .A2(_06463_),
    .B1(_06497_),
    .C1(_06810_),
    .X(_06841_));
 sky130_fd_sc_hd__nand2_4 _12403_ (.A(_06840_),
    .B(_06841_),
    .Y(\CPU_result_a3[4] ));
 sky130_fd_sc_hd__o22a_4 _12404_ (.A1(\CPU_dmem_rd_data_a5[4] ),
    .A2(CPU_valid_a3),
    .B1(_06173_),
    .B2(\CPU_result_a3[4] ),
    .X(_06842_));
 sky130_fd_sc_hd__inv_2 _12405_ (.A(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__buf_2 _12406_ (.A(_06628_),
    .X(_06844_));
 sky130_fd_sc_hd__nor2_4 _12407_ (.A(\CPU_Xreg_value_a4[1][4] ),
    .B(_06544_),
    .Y(_06845_));
 sky130_fd_sc_hd__a211o_4 _12408_ (.A1(_06783_),
    .A2(_06843_),
    .B1(_06844_),
    .C1(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__inv_2 _12409_ (.A(_06846_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_4 _12410_ (.A(_06278_),
    .B(_06279_),
    .Y(_06847_));
 sky130_fd_sc_hd__a21o_4 _12411_ (.A1(\CPU_src2_value_a3[3] ),
    .A2(\CPU_src1_value_a3[3] ),
    .B1(_06465_),
    .X(_06848_));
 sky130_fd_sc_hd__nand2_4 _12412_ (.A(_06475_),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__o21a_4 _12413_ (.A1(_06475_),
    .A2(_06848_),
    .B1(_06499_),
    .X(_06850_));
 sky130_fd_sc_hd__a32o_4 _12414_ (.A1(_06280_),
    .A2(_06180_),
    .A3(_06847_),
    .B1(_06849_),
    .B2(_06850_),
    .X(\CPU_result_a3[3] ));
 sky130_fd_sc_hd__o22a_4 _12415_ (.A1(\CPU_dmem_rd_data_a5[3] ),
    .A2(CPU_valid_a3),
    .B1(_06173_),
    .B2(\CPU_result_a3[3] ),
    .X(_06851_));
 sky130_fd_sc_hd__inv_2 _12416_ (.A(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__nor2_4 _12417_ (.A(\CPU_Xreg_value_a4[1][3] ),
    .B(_06544_),
    .Y(_06853_));
 sky130_fd_sc_hd__a211o_4 _12418_ (.A1(_06504_),
    .A2(_06852_),
    .B1(_06844_),
    .C1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__inv_2 _12419_ (.A(_06854_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_4 _12420_ (.A(_06275_),
    .B(_06276_),
    .Y(_06855_));
 sky130_fd_sc_hd__a21o_4 _12421_ (.A1(\CPU_src2_value_a3[2] ),
    .A2(\CPU_src1_value_a3[2] ),
    .B1(_06467_),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_4 _12422_ (.A(_06474_),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__o21a_4 _12423_ (.A1(_06474_),
    .A2(_06856_),
    .B1(_06499_),
    .X(_06858_));
 sky130_fd_sc_hd__a32o_4 _12424_ (.A1(_06277_),
    .A2(_06180_),
    .A3(_06855_),
    .B1(_06857_),
    .B2(_06858_),
    .X(\CPU_result_a3[2] ));
 sky130_fd_sc_hd__o22a_4 _12425_ (.A1(\CPU_dmem_rd_data_a5[2] ),
    .A2(CPU_valid_a3),
    .B1(_06173_),
    .B2(\CPU_result_a3[2] ),
    .X(_06859_));
 sky130_fd_sc_hd__inv_2 _12426_ (.A(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__nor2_4 _12427_ (.A(\CPU_Xreg_value_a4[1][2] ),
    .B(_06544_),
    .Y(_06861_));
 sky130_fd_sc_hd__a211o_4 _12428_ (.A1(_06504_),
    .A2(_06860_),
    .B1(_06844_),
    .C1(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__inv_2 _12429_ (.A(_06862_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_4 _12430_ (.A(_06470_),
    .B(_06472_),
    .Y(_06863_));
 sky130_fd_sc_hd__o21ai_4 _12431_ (.A1(_06271_),
    .A2(_06272_),
    .B1(_06273_),
    .Y(_06864_));
 sky130_fd_sc_hd__and2_4 _12432_ (.A(_06274_),
    .B(_06581_),
    .X(_06865_));
 sky130_fd_sc_hd__a32o_4 _12433_ (.A1(_06473_),
    .A2(_06577_),
    .A3(_06863_),
    .B1(_06864_),
    .B2(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__o22a_4 _12434_ (.A1(\CPU_dmem_rd_data_a5[1] ),
    .A2(_06171_),
    .B1(_06173_),
    .B2(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__inv_2 _12435_ (.A(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__nor2_4 _12436_ (.A(\CPU_Xreg_value_a4[1][1] ),
    .B(_06544_),
    .Y(_06869_));
 sky130_fd_sc_hd__a211o_4 _12437_ (.A1(_06504_),
    .A2(_06868_),
    .B1(_06844_),
    .C1(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__inv_2 _12438_ (.A(_06870_),
    .Y(_00975_));
 sky130_fd_sc_hd__and2_4 _12439_ (.A(_06271_),
    .B(\CPU_imm_a3[0] ),
    .X(_06871_));
 sky130_fd_sc_hd__a21oi_4 _12440_ (.A1(\CPU_src1_value_a3[0] ),
    .A2(_06272_),
    .B1(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__inv_2 _12441_ (.A(_06470_),
    .Y(_06873_));
 sky130_fd_sc_hd__a211o_4 _12442_ (.A1(_06469_),
    .A2(_06271_),
    .B1(_06495_),
    .C1(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__inv_2 _12443_ (.A(CPU_is_slti_a3),
    .Y(_06875_));
 sky130_fd_sc_hd__a211o_4 _12444_ (.A1(_06468_),
    .A2(\CPU_src1_value_a3[1] ),
    .B1(_06469_),
    .C1(\CPU_src1_value_a3[0] ),
    .X(_06876_));
 sky130_fd_sc_hd__a32o_4 _12445_ (.A1(_06471_),
    .A2(_06856_),
    .A3(_06876_),
    .B1(_06466_),
    .B2(\CPU_src1_value_a3[2] ),
    .X(_06877_));
 sky130_fd_sc_hd__a22oi_4 _12446_ (.A1(_06464_),
    .A2(\CPU_src1_value_a3[3] ),
    .B1(_06848_),
    .B2(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__and4_4 _12447_ (.A(_06456_),
    .B(_06462_),
    .C(_06458_),
    .D(_06463_),
    .X(_06879_));
 sky130_fd_sc_hd__inv_2 _12448_ (.A(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__or3_4 _12449_ (.A(_06294_),
    .B(\CPU_src2_value_a3[4] ),
    .C(_06832_),
    .X(_06881_));
 sky130_fd_sc_hd__o22a_4 _12450_ (.A1(\CPU_src2_value_a3[6] ),
    .A2(_06285_),
    .B1(\CPU_src2_value_a3[5] ),
    .B2(_06288_),
    .X(_06882_));
 sky130_fd_sc_hd__and2_4 _12451_ (.A(_06881_),
    .B(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__o32a_4 _12452_ (.A1(_06455_),
    .A2(_06457_),
    .A3(_06883_),
    .B1(\CPU_src2_value_a3[7] ),
    .B2(_06282_),
    .X(_06884_));
 sky130_fd_sc_hd__o21a_4 _12453_ (.A1(_06878_),
    .A2(_06880_),
    .B1(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__inv_2 _12454_ (.A(_06442_),
    .Y(_06886_));
 sky130_fd_sc_hd__inv_2 _12455_ (.A(_06443_),
    .Y(_06887_));
 sky130_fd_sc_hd__or2_4 _12456_ (.A(_06430_),
    .B(_06433_),
    .X(_06888_));
 sky130_fd_sc_hd__or4_4 _12457_ (.A(_06432_),
    .B(_06886_),
    .C(_06887_),
    .D(_06888_),
    .X(_06889_));
 sky130_fd_sc_hd__inv_2 _12458_ (.A(\CPU_src1_value_a3[11] ),
    .Y(_06890_));
 sky130_fd_sc_hd__and3_4 _12459_ (.A(\CPU_src1_value_a3[8] ),
    .B(_06437_),
    .C(_06443_),
    .X(_06891_));
 sky130_fd_sc_hd__a211o_4 _12460_ (.A1(_06435_),
    .A2(\CPU_src1_value_a3[9] ),
    .B1(_06432_),
    .C1(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__inv_2 _12461_ (.A(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__o22a_4 _12462_ (.A1(\CPU_src2_value_a3[11] ),
    .A2(_06890_),
    .B1(_06888_),
    .B2(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__o21a_4 _12463_ (.A1(_06885_),
    .A2(_06889_),
    .B1(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__inv_2 _12464_ (.A(_06422_),
    .Y(_06896_));
 sky130_fd_sc_hd__inv_2 _12465_ (.A(_06423_),
    .Y(_06897_));
 sky130_fd_sc_hd__inv_2 _12466_ (.A(_06410_),
    .Y(_06898_));
 sky130_fd_sc_hd__or2_4 _12467_ (.A(_06898_),
    .B(_06413_),
    .X(_06899_));
 sky130_fd_sc_hd__or4_4 _12468_ (.A(_06412_),
    .B(_06896_),
    .C(_06897_),
    .D(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__and3_4 _12469_ (.A(\CPU_src1_value_a3[12] ),
    .B(_06417_),
    .C(_06423_),
    .X(_06901_));
 sky130_fd_sc_hd__a211o_4 _12470_ (.A1(_06415_),
    .A2(\CPU_src1_value_a3[13] ),
    .B1(_06412_),
    .C1(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__inv_2 _12471_ (.A(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__o22a_4 _12472_ (.A1(\CPU_src2_value_a3[15] ),
    .A2(_06233_),
    .B1(_06899_),
    .B2(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__o21ai_4 _12473_ (.A1(_06895_),
    .A2(_06900_),
    .B1(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__and4_4 _12474_ (.A(_06346_),
    .B(_06353_),
    .C(_06354_),
    .D(_06493_),
    .X(_06906_));
 sky130_fd_sc_hd__and4_4 _12475_ (.A(_06406_),
    .B(_06407_),
    .C(_06396_),
    .D(_06398_),
    .X(_06907_));
 sky130_fd_sc_hd__and4_4 _12476_ (.A(_06367_),
    .B(_06369_),
    .C(_06373_),
    .D(_06374_),
    .X(_06908_));
 sky130_fd_sc_hd__and4_4 _12477_ (.A(_06387_),
    .B(_06388_),
    .C(_06376_),
    .D(_06379_),
    .X(_06909_));
 sky130_fd_sc_hd__and4_4 _12478_ (.A(_06906_),
    .B(_06907_),
    .C(_06908_),
    .D(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__or3_4 _12479_ (.A(_06200_),
    .B(\CPU_src2_value_a3[28] ),
    .C(_06352_),
    .X(_06911_));
 sky130_fd_sc_hd__o22a_4 _12480_ (.A1(\CPU_src2_value_a3[30] ),
    .A2(_06181_),
    .B1(\CPU_src2_value_a3[29] ),
    .B2(_06197_),
    .X(_06912_));
 sky130_fd_sc_hd__a211o_4 _12481_ (.A1(_06911_),
    .A2(_06912_),
    .B1(_06345_),
    .C1(_06491_),
    .X(_06913_));
 sky130_fd_sc_hd__inv_2 _12482_ (.A(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__and2_4 _12483_ (.A(_06399_),
    .B(\CPU_src1_value_a3[17] ),
    .X(_06915_));
 sky130_fd_sc_hd__and3_4 _12484_ (.A(\CPU_src1_value_a3[16] ),
    .B(_06401_),
    .C(_06407_),
    .X(_06916_));
 sky130_fd_sc_hd__a211o_4 _12485_ (.A1(_06392_),
    .A2(\CPU_src1_value_a3[18] ),
    .B1(_06915_),
    .C1(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__a32o_4 _12486_ (.A1(_06396_),
    .A2(_06397_),
    .A3(_06917_),
    .B1(_06390_),
    .B2(\CPU_src1_value_a3[19] ),
    .X(_06918_));
 sky130_fd_sc_hd__nor2_4 _12487_ (.A(\CPU_src2_value_a3[23] ),
    .B(_06221_),
    .Y(_06919_));
 sky130_fd_sc_hd__inv_2 _12488_ (.A(_06388_),
    .Y(_06920_));
 sky130_fd_sc_hd__or3_4 _12489_ (.A(_06218_),
    .B(\CPU_src2_value_a3[20] ),
    .C(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__o22a_4 _12490_ (.A1(\CPU_src2_value_a3[22] ),
    .A2(_06312_),
    .B1(\CPU_src2_value_a3[21] ),
    .B2(_06216_),
    .X(_06922_));
 sky130_fd_sc_hd__inv_2 _12491_ (.A(_06376_),
    .Y(_06923_));
 sky130_fd_sc_hd__a211o_4 _12492_ (.A1(_06921_),
    .A2(_06922_),
    .B1(_06923_),
    .C1(_06378_),
    .X(_06924_));
 sky130_fd_sc_hd__inv_2 _12493_ (.A(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__a211o_4 _12494_ (.A1(_06909_),
    .A2(_06918_),
    .B1(_06919_),
    .C1(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__or3_4 _12495_ (.A(_06205_),
    .B(\CPU_src2_value_a3[24] ),
    .C(_06579_),
    .X(_06927_));
 sky130_fd_sc_hd__o22a_4 _12496_ (.A1(\CPU_src2_value_a3[26] ),
    .A2(_06211_),
    .B1(\CPU_src2_value_a3[25] ),
    .B2(_06204_),
    .X(_06928_));
 sky130_fd_sc_hd__a211o_4 _12497_ (.A1(_06927_),
    .A2(_06928_),
    .B1(_06366_),
    .C1(_06368_),
    .X(_06929_));
 sky130_fd_sc_hd__inv_2 _12498_ (.A(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__and2_4 _12499_ (.A(_06355_),
    .B(\CPU_src1_value_a3[27] ),
    .X(_06931_));
 sky130_fd_sc_hd__a211o_4 _12500_ (.A1(_06908_),
    .A2(_06926_),
    .B1(_06930_),
    .C1(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__and2_4 _12501_ (.A(_06906_),
    .B(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__a2111o_4 _12502_ (.A1(_06905_),
    .A2(_06910_),
    .B1(_06490_),
    .C1(_06914_),
    .D1(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__or2_4 _12503_ (.A(_06492_),
    .B(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__and4_4 _12504_ (.A(_06875_),
    .B(CPU_is_slt_a3),
    .C(_06489_),
    .D(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__and2_4 _12505_ (.A(\CPU_src1_value_a3[7] ),
    .B(\CPU_src1_value_a3[6] ),
    .X(_06937_));
 sky130_fd_sc_hd__or2_4 _12506_ (.A(_06283_),
    .B(_06286_),
    .X(_06938_));
 sky130_fd_sc_hd__o21a_4 _12507_ (.A1(_06271_),
    .A2(\CPU_imm_a3[0] ),
    .B1(_06273_),
    .X(_06939_));
 sky130_fd_sc_hd__a2bb2o_4 _12508_ (.A1_N(\CPU_src1_value_a3[1] ),
    .A2_N(_06270_),
    .B1(_06267_),
    .B2(\CPU_imm_a3[2] ),
    .X(_06940_));
 sky130_fd_sc_hd__o22a_4 _12509_ (.A1(_06267_),
    .A2(\CPU_imm_a3[2] ),
    .B1(_06265_),
    .B2(\CPU_imm_a3[3] ),
    .X(_06941_));
 sky130_fd_sc_hd__o21a_4 _12510_ (.A1(_06939_),
    .A2(_06940_),
    .B1(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__a211o_4 _12511_ (.A1(_06265_),
    .A2(\CPU_imm_a3[3] ),
    .B1(_06295_),
    .C1(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__a32o_4 _12512_ (.A1(_06293_),
    .A2(_06296_),
    .A3(_06943_),
    .B1(_06288_),
    .B2(_06194_),
    .X(_06944_));
 sky130_fd_sc_hd__inv_2 _12513_ (.A(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__o22a_4 _12514_ (.A1(_06187_),
    .A2(_06937_),
    .B1(_06938_),
    .B2(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__inv_2 _12515_ (.A(_06247_),
    .Y(_06947_));
 sky130_fd_sc_hd__or4_4 _12516_ (.A(_06947_),
    .B(_06249_),
    .C(_06260_),
    .D(_06262_),
    .X(_06948_));
 sky130_fd_sc_hd__or3_4 _12517_ (.A(_06248_),
    .B(_06253_),
    .C(_06260_),
    .X(_06949_));
 sky130_fd_sc_hd__a32o_4 _12518_ (.A1(_06195_),
    .A2(_06247_),
    .A3(_06949_),
    .B1(_06890_),
    .B2(\CPU_imm_a3[11] ),
    .X(_06950_));
 sky130_fd_sc_hd__inv_2 _12519_ (.A(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__o21a_4 _12520_ (.A1(_06946_),
    .A2(_06948_),
    .B1(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__or4_4 _12521_ (.A(_06235_),
    .B(_06239_),
    .C(_06237_),
    .D(_06242_),
    .X(_06953_));
 sky130_fd_sc_hd__and4_4 _12522_ (.A(_06236_),
    .B(_06240_),
    .C(\CPU_src1_value_a3[14] ),
    .D(\CPU_src1_value_a3[12] ),
    .X(_06954_));
 sky130_fd_sc_hd__o22a_4 _12523_ (.A1(_06952_),
    .A2(_06953_),
    .B1(_06188_),
    .B2(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__or4_4 _12524_ (.A(_06316_),
    .B(_06313_),
    .C(_06657_),
    .D(_06655_),
    .X(_06956_));
 sky130_fd_sc_hd__nand2_4 _12525_ (.A(_06583_),
    .B(_06212_),
    .Y(_06957_));
 sky130_fd_sc_hd__or3_4 _12526_ (.A(_06547_),
    .B(_06198_),
    .C(_06213_),
    .X(_06958_));
 sky130_fd_sc_hd__or4_4 _12527_ (.A(_06315_),
    .B(_06310_),
    .C(_06656_),
    .D(_06654_),
    .X(_06959_));
 sky130_fd_sc_hd__or4_4 _12528_ (.A(_06340_),
    .B(_06957_),
    .C(_06958_),
    .D(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__or4_4 _12529_ (.A(_06196_),
    .B(_06201_),
    .C(_06956_),
    .D(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__or4_4 _12530_ (.A(_06199_),
    .B(_06211_),
    .C(_06206_),
    .D(_06312_),
    .X(_06962_));
 sky130_fd_sc_hd__or3_4 _12531_ (.A(_06218_),
    .B(_06324_),
    .C(_06320_),
    .X(_06963_));
 sky130_fd_sc_hd__or4_4 _12532_ (.A(_06338_),
    .B(_06181_),
    .C(_06962_),
    .D(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__or3_4 _12533_ (.A(_06958_),
    .B(_06964_),
    .C(_06959_),
    .X(_06965_));
 sky130_fd_sc_hd__a2bb2o_4 _12534_ (.A1_N(_06955_),
    .A2_N(_06961_),
    .B1(_06195_),
    .B2(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__inv_2 _12535_ (.A(_06276_),
    .Y(_06967_));
 sky130_fd_sc_hd__inv_2 _12536_ (.A(_06279_),
    .Y(_06968_));
 sky130_fd_sc_hd__or4_4 _12537_ (.A(_06295_),
    .B(_06871_),
    .C(_06967_),
    .D(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__inv_2 _12538_ (.A(_06939_),
    .Y(_06970_));
 sky130_fd_sc_hd__or4_4 _12539_ (.A(_06834_),
    .B(_06297_),
    .C(_06938_),
    .D(_06970_),
    .X(_06971_));
 sky130_fd_sc_hd__or4_4 _12540_ (.A(_06948_),
    .B(_06969_),
    .C(_06953_),
    .D(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__o22a_4 _12541_ (.A1(\CPU_src1_value_a3[31] ),
    .A2(_06189_),
    .B1(_06961_),
    .B2(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__and2_4 _12542_ (.A(_06966_),
    .B(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__or3_4 _12543_ (.A(_06875_),
    .B(_06339_),
    .C(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__inv_2 _12544_ (.A(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__or3_4 _12545_ (.A(CPU_is_add_a3),
    .B(_06936_),
    .C(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__and3_4 _12546_ (.A(_06174_),
    .B(_06874_),
    .C(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__a21oi_4 _12547_ (.A1(_06582_),
    .A2(_06872_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__o22a_4 _12548_ (.A1(\CPU_dmem_rd_data_a5[0] ),
    .A2(CPU_valid_a3),
    .B1(_06173_),
    .B2(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__buf_2 _12549_ (.A(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__inv_2 _12550_ (.A(\CPU_Xreg_value_a4[1][0] ),
    .Y(_06982_));
 sky130_fd_sc_hd__nor2_4 _12551_ (.A(_06982_),
    .B(_06169_),
    .Y(_06983_));
 sky130_fd_sc_hd__a211o_4 _12552_ (.A1(_06169_),
    .A2(_06981_),
    .B1(_06140_),
    .C1(_06983_),
    .X(_00974_));
 sky130_fd_sc_hd__buf_2 _12553_ (.A(_06503_),
    .X(_06984_));
 sky130_fd_sc_hd__inv_2 _12554_ (.A(_06151_),
    .Y(_06985_));
 sky130_fd_sc_hd__or2_4 _12555_ (.A(_06149_),
    .B(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__or2_4 _12556_ (.A(_06148_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__nor2_4 _12557_ (.A(_06166_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__buf_2 _12558_ (.A(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__buf_2 _12559_ (.A(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__buf_2 _12560_ (.A(_06989_),
    .X(_06991_));
 sky130_fd_sc_hd__nor2_4 _12561_ (.A(\CPU_Xreg_value_a4[2][31] ),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__a211o_4 _12562_ (.A1(_06984_),
    .A2(_06990_),
    .B1(_06844_),
    .C1(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__inv_2 _12563_ (.A(_06993_),
    .Y(_00973_));
 sky130_fd_sc_hd__buf_2 _12564_ (.A(_06515_),
    .X(_06994_));
 sky130_fd_sc_hd__nor2_4 _12565_ (.A(\CPU_Xreg_value_a4[2][30] ),
    .B(_06991_),
    .Y(_06995_));
 sky130_fd_sc_hd__a211o_4 _12566_ (.A1(_06994_),
    .A2(_06990_),
    .B1(_06844_),
    .C1(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__inv_2 _12567_ (.A(_06996_),
    .Y(_00972_));
 sky130_fd_sc_hd__buf_2 _12568_ (.A(_06531_),
    .X(_06997_));
 sky130_fd_sc_hd__buf_2 _12569_ (.A(_06628_),
    .X(_06998_));
 sky130_fd_sc_hd__nor2_4 _12570_ (.A(\CPU_Xreg_value_a4[2][29] ),
    .B(_06991_),
    .Y(_06999_));
 sky130_fd_sc_hd__a211o_4 _12571_ (.A1(_06997_),
    .A2(_06990_),
    .B1(_06998_),
    .C1(_06999_),
    .X(_07000_));
 sky130_fd_sc_hd__inv_2 _12572_ (.A(_07000_),
    .Y(_00971_));
 sky130_fd_sc_hd__buf_2 _12573_ (.A(_06539_),
    .X(_07001_));
 sky130_fd_sc_hd__buf_2 _12574_ (.A(_06989_),
    .X(_07002_));
 sky130_fd_sc_hd__nor2_4 _12575_ (.A(\CPU_Xreg_value_a4[2][28] ),
    .B(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__a211o_4 _12576_ (.A1(_07001_),
    .A2(_06990_),
    .B1(_06998_),
    .C1(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__inv_2 _12577_ (.A(_07004_),
    .Y(_00970_));
 sky130_fd_sc_hd__buf_2 _12578_ (.A(_06564_),
    .X(_07005_));
 sky130_fd_sc_hd__buf_2 _12579_ (.A(_06988_),
    .X(_07006_));
 sky130_fd_sc_hd__buf_2 _12580_ (.A(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__nor2_4 _12581_ (.A(\CPU_Xreg_value_a4[2][27] ),
    .B(_07002_),
    .Y(_07008_));
 sky130_fd_sc_hd__a211o_4 _12582_ (.A1(_07005_),
    .A2(_07007_),
    .B1(_06998_),
    .C1(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__inv_2 _12583_ (.A(_07009_),
    .Y(_00969_));
 sky130_fd_sc_hd__buf_2 _12584_ (.A(_06574_),
    .X(_07010_));
 sky130_fd_sc_hd__nor2_4 _12585_ (.A(\CPU_Xreg_value_a4[2][26] ),
    .B(_07002_),
    .Y(_07011_));
 sky130_fd_sc_hd__a211o_4 _12586_ (.A1(_07010_),
    .A2(_07007_),
    .B1(_06998_),
    .C1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__inv_2 _12587_ (.A(_07012_),
    .Y(_00968_));
 sky130_fd_sc_hd__buf_2 _12588_ (.A(_06589_),
    .X(_07013_));
 sky130_fd_sc_hd__nor2_4 _12589_ (.A(\CPU_Xreg_value_a4[2][25] ),
    .B(_07002_),
    .Y(_07014_));
 sky130_fd_sc_hd__a211o_4 _12590_ (.A1(_07013_),
    .A2(_07007_),
    .B1(_06998_),
    .C1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__inv_2 _12591_ (.A(_07015_),
    .Y(_00967_));
 sky130_fd_sc_hd__buf_2 _12592_ (.A(_06599_),
    .X(_07016_));
 sky130_fd_sc_hd__nor2_4 _12593_ (.A(\CPU_Xreg_value_a4[2][24] ),
    .B(_07002_),
    .Y(_07017_));
 sky130_fd_sc_hd__a211o_4 _12594_ (.A1(_07016_),
    .A2(_07007_),
    .B1(_06998_),
    .C1(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__inv_2 _12595_ (.A(_07018_),
    .Y(_00966_));
 sky130_fd_sc_hd__buf_2 _12596_ (.A(_06619_),
    .X(_07019_));
 sky130_fd_sc_hd__buf_2 _12597_ (.A(_06628_),
    .X(_07020_));
 sky130_fd_sc_hd__nor2_4 _12598_ (.A(\CPU_Xreg_value_a4[2][23] ),
    .B(_07002_),
    .Y(_07021_));
 sky130_fd_sc_hd__a211o_4 _12599_ (.A1(_07019_),
    .A2(_07007_),
    .B1(_07020_),
    .C1(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__inv_2 _12600_ (.A(_07022_),
    .Y(_00965_));
 sky130_fd_sc_hd__buf_2 _12601_ (.A(_06627_),
    .X(_07023_));
 sky130_fd_sc_hd__buf_2 _12602_ (.A(_06989_),
    .X(_07024_));
 sky130_fd_sc_hd__nor2_4 _12603_ (.A(\CPU_Xreg_value_a4[2][22] ),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__a211o_4 _12604_ (.A1(_07023_),
    .A2(_07007_),
    .B1(_07020_),
    .C1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__inv_2 _12605_ (.A(_07026_),
    .Y(_00964_));
 sky130_fd_sc_hd__buf_2 _12606_ (.A(_06642_),
    .X(_07027_));
 sky130_fd_sc_hd__buf_2 _12607_ (.A(_07006_),
    .X(_07028_));
 sky130_fd_sc_hd__nor2_4 _12608_ (.A(\CPU_Xreg_value_a4[2][21] ),
    .B(_07024_),
    .Y(_07029_));
 sky130_fd_sc_hd__a211o_4 _12609_ (.A1(_07027_),
    .A2(_07028_),
    .B1(_07020_),
    .C1(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__inv_2 _12610_ (.A(_07030_),
    .Y(_00963_));
 sky130_fd_sc_hd__buf_2 _12611_ (.A(_06651_),
    .X(_07031_));
 sky130_fd_sc_hd__nor2_4 _12612_ (.A(\CPU_Xreg_value_a4[2][20] ),
    .B(_07024_),
    .Y(_07032_));
 sky130_fd_sc_hd__a211o_4 _12613_ (.A1(_07031_),
    .A2(_07028_),
    .B1(_07020_),
    .C1(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__inv_2 _12614_ (.A(_07033_),
    .Y(_00962_));
 sky130_fd_sc_hd__buf_2 _12615_ (.A(_06673_),
    .X(_07034_));
 sky130_fd_sc_hd__nor2_4 _12616_ (.A(\CPU_Xreg_value_a4[2][19] ),
    .B(_07024_),
    .Y(_07035_));
 sky130_fd_sc_hd__a211o_4 _12617_ (.A1(_07034_),
    .A2(_07028_),
    .B1(_07020_),
    .C1(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__inv_2 _12618_ (.A(_07036_),
    .Y(_00961_));
 sky130_fd_sc_hd__buf_2 _12619_ (.A(_06682_),
    .X(_07037_));
 sky130_fd_sc_hd__nor2_4 _12620_ (.A(\CPU_Xreg_value_a4[2][18] ),
    .B(_07024_),
    .Y(_07038_));
 sky130_fd_sc_hd__a211o_4 _12621_ (.A1(_07037_),
    .A2(_07028_),
    .B1(_07020_),
    .C1(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__inv_2 _12622_ (.A(_07039_),
    .Y(_00960_));
 sky130_fd_sc_hd__buf_2 _12623_ (.A(_06692_),
    .X(_07040_));
 sky130_fd_sc_hd__buf_2 _12624_ (.A(_06101_),
    .X(_07041_));
 sky130_fd_sc_hd__buf_2 _12625_ (.A(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__nor2_4 _12626_ (.A(\CPU_Xreg_value_a4[2][17] ),
    .B(_07024_),
    .Y(_07043_));
 sky130_fd_sc_hd__a211o_4 _12627_ (.A1(_07040_),
    .A2(_07028_),
    .B1(_07042_),
    .C1(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__inv_2 _12628_ (.A(_07044_),
    .Y(_00959_));
 sky130_fd_sc_hd__buf_2 _12629_ (.A(_06701_),
    .X(_07045_));
 sky130_fd_sc_hd__buf_2 _12630_ (.A(_06988_),
    .X(_07046_));
 sky130_fd_sc_hd__nor2_4 _12631_ (.A(\CPU_Xreg_value_a4[2][16] ),
    .B(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__a211o_4 _12632_ (.A1(_07045_),
    .A2(_07028_),
    .B1(_07042_),
    .C1(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__inv_2 _12633_ (.A(_07048_),
    .Y(_00958_));
 sky130_fd_sc_hd__buf_2 _12634_ (.A(_06724_),
    .X(_07049_));
 sky130_fd_sc_hd__buf_2 _12635_ (.A(_06989_),
    .X(_07050_));
 sky130_fd_sc_hd__nor2_4 _12636_ (.A(\CPU_Xreg_value_a4[2][15] ),
    .B(_07046_),
    .Y(_07051_));
 sky130_fd_sc_hd__a211o_4 _12637_ (.A1(_07049_),
    .A2(_07050_),
    .B1(_07042_),
    .C1(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__inv_2 _12638_ (.A(_07052_),
    .Y(_00957_));
 sky130_fd_sc_hd__buf_2 _12639_ (.A(_06733_),
    .X(_07053_));
 sky130_fd_sc_hd__nor2_4 _12640_ (.A(\CPU_Xreg_value_a4[2][14] ),
    .B(_07046_),
    .Y(_07054_));
 sky130_fd_sc_hd__a211o_4 _12641_ (.A1(_07053_),
    .A2(_07050_),
    .B1(_07042_),
    .C1(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__inv_2 _12642_ (.A(_07055_),
    .Y(_00956_));
 sky130_fd_sc_hd__buf_2 _12643_ (.A(_06743_),
    .X(_07056_));
 sky130_fd_sc_hd__nor2_4 _12644_ (.A(\CPU_Xreg_value_a4[2][13] ),
    .B(_07046_),
    .Y(_07057_));
 sky130_fd_sc_hd__a211o_4 _12645_ (.A1(_07056_),
    .A2(_07050_),
    .B1(_07042_),
    .C1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__inv_2 _12646_ (.A(_07058_),
    .Y(_00955_));
 sky130_fd_sc_hd__buf_2 _12647_ (.A(_06752_),
    .X(_07059_));
 sky130_fd_sc_hd__nor2_4 _12648_ (.A(\CPU_Xreg_value_a4[2][12] ),
    .B(_07046_),
    .Y(_07060_));
 sky130_fd_sc_hd__a211o_4 _12649_ (.A1(_07059_),
    .A2(_07050_),
    .B1(_07042_),
    .C1(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__inv_2 _12650_ (.A(_07061_),
    .Y(_00954_));
 sky130_fd_sc_hd__buf_2 _12651_ (.A(_06770_),
    .X(_07062_));
 sky130_fd_sc_hd__buf_2 _12652_ (.A(_07041_),
    .X(_07063_));
 sky130_fd_sc_hd__nor2_4 _12653_ (.A(\CPU_Xreg_value_a4[2][11] ),
    .B(_07046_),
    .Y(_07064_));
 sky130_fd_sc_hd__a211o_4 _12654_ (.A1(_07062_),
    .A2(_07050_),
    .B1(_07063_),
    .C1(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__inv_2 _12655_ (.A(_07065_),
    .Y(_00953_));
 sky130_fd_sc_hd__buf_2 _12656_ (.A(_06778_),
    .X(_07066_));
 sky130_fd_sc_hd__buf_2 _12657_ (.A(_06988_),
    .X(_07067_));
 sky130_fd_sc_hd__nor2_4 _12658_ (.A(\CPU_Xreg_value_a4[2][10] ),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a211o_4 _12659_ (.A1(_07066_),
    .A2(_07050_),
    .B1(_07063_),
    .C1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__inv_2 _12660_ (.A(_07069_),
    .Y(_00952_));
 sky130_fd_sc_hd__buf_2 _12661_ (.A(_06791_),
    .X(_07070_));
 sky130_fd_sc_hd__buf_2 _12662_ (.A(_06989_),
    .X(_07071_));
 sky130_fd_sc_hd__nor2_4 _12663_ (.A(\CPU_Xreg_value_a4[2][9] ),
    .B(_07067_),
    .Y(_07072_));
 sky130_fd_sc_hd__a211o_4 _12664_ (.A1(_07070_),
    .A2(_07071_),
    .B1(_07063_),
    .C1(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__inv_2 _12665_ (.A(_07073_),
    .Y(_00951_));
 sky130_fd_sc_hd__buf_2 _12666_ (.A(_06799_),
    .X(_07074_));
 sky130_fd_sc_hd__nor2_4 _12667_ (.A(\CPU_Xreg_value_a4[2][8] ),
    .B(_07067_),
    .Y(_07075_));
 sky130_fd_sc_hd__a211o_4 _12668_ (.A1(_07074_),
    .A2(_07071_),
    .B1(_07063_),
    .C1(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__inv_2 _12669_ (.A(_07076_),
    .Y(_00950_));
 sky130_fd_sc_hd__buf_2 _12670_ (.A(_06820_),
    .X(_07077_));
 sky130_fd_sc_hd__nor2_4 _12671_ (.A(\CPU_Xreg_value_a4[2][7] ),
    .B(_07067_),
    .Y(_07078_));
 sky130_fd_sc_hd__a211o_4 _12672_ (.A1(_07077_),
    .A2(_07071_),
    .B1(_07063_),
    .C1(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__inv_2 _12673_ (.A(_07079_),
    .Y(_00949_));
 sky130_fd_sc_hd__buf_2 _12674_ (.A(_06828_),
    .X(_07080_));
 sky130_fd_sc_hd__nor2_4 _12675_ (.A(\CPU_Xreg_value_a4[2][6] ),
    .B(_07067_),
    .Y(_07081_));
 sky130_fd_sc_hd__a211o_4 _12676_ (.A1(_07080_),
    .A2(_07071_),
    .B1(_07063_),
    .C1(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__inv_2 _12677_ (.A(_07082_),
    .Y(_00948_));
 sky130_fd_sc_hd__buf_2 _12678_ (.A(_06837_),
    .X(_07083_));
 sky130_fd_sc_hd__buf_2 _12679_ (.A(_07041_),
    .X(_07084_));
 sky130_fd_sc_hd__nor2_4 _12680_ (.A(\CPU_Xreg_value_a4[2][5] ),
    .B(_07067_),
    .Y(_07085_));
 sky130_fd_sc_hd__a211o_4 _12681_ (.A1(_07083_),
    .A2(_07071_),
    .B1(_07084_),
    .C1(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__inv_2 _12682_ (.A(_07086_),
    .Y(_00947_));
 sky130_fd_sc_hd__buf_2 _12683_ (.A(_06843_),
    .X(_07087_));
 sky130_fd_sc_hd__nor2_4 _12684_ (.A(\CPU_Xreg_value_a4[2][4] ),
    .B(_07006_),
    .Y(_07088_));
 sky130_fd_sc_hd__a211o_4 _12685_ (.A1(_07087_),
    .A2(_07071_),
    .B1(_07084_),
    .C1(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__inv_2 _12686_ (.A(_07089_),
    .Y(_00946_));
 sky130_fd_sc_hd__buf_2 _12687_ (.A(_06852_),
    .X(_07090_));
 sky130_fd_sc_hd__nor2_4 _12688_ (.A(\CPU_Xreg_value_a4[2][3] ),
    .B(_07006_),
    .Y(_07091_));
 sky130_fd_sc_hd__a211o_4 _12689_ (.A1(_07090_),
    .A2(_06991_),
    .B1(_07084_),
    .C1(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__inv_2 _12690_ (.A(_07092_),
    .Y(_00945_));
 sky130_fd_sc_hd__buf_2 _12691_ (.A(_06860_),
    .X(_07093_));
 sky130_fd_sc_hd__nor2_4 _12692_ (.A(\CPU_Xreg_value_a4[2][2] ),
    .B(_07006_),
    .Y(_07094_));
 sky130_fd_sc_hd__a211o_4 _12693_ (.A1(_07093_),
    .A2(_06991_),
    .B1(_07084_),
    .C1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__inv_2 _12694_ (.A(_07095_),
    .Y(_00944_));
 sky130_fd_sc_hd__buf_2 _12695_ (.A(_06867_),
    .X(_07096_));
 sky130_fd_sc_hd__buf_2 _12696_ (.A(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__inv_2 _12697_ (.A(\CPU_Xreg_value_a4[2][1] ),
    .Y(_07098_));
 sky130_fd_sc_hd__nor2_4 _12698_ (.A(_07098_),
    .B(_06990_),
    .Y(_07099_));
 sky130_fd_sc_hd__a211o_4 _12699_ (.A1(_07097_),
    .A2(_06990_),
    .B1(_06140_),
    .C1(_07099_),
    .X(_00943_));
 sky130_fd_sc_hd__inv_2 _12700_ (.A(_06980_),
    .Y(_07100_));
 sky130_fd_sc_hd__buf_2 _12701_ (.A(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__nor2_4 _12702_ (.A(\CPU_Xreg_value_a4[2][0] ),
    .B(_07006_),
    .Y(_07102_));
 sky130_fd_sc_hd__a211o_4 _12703_ (.A1(_07101_),
    .A2(_06991_),
    .B1(_07084_),
    .C1(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__inv_2 _12704_ (.A(_07103_),
    .Y(_00942_));
 sky130_fd_sc_hd__or2_4 _12705_ (.A(_06150_),
    .B(_06985_),
    .X(_07104_));
 sky130_fd_sc_hd__or2_4 _12706_ (.A(_06148_),
    .B(_07104_),
    .X(_07105_));
 sky130_fd_sc_hd__nor2_4 _12707_ (.A(_06166_),
    .B(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__buf_2 _12708_ (.A(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__buf_2 _12709_ (.A(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__buf_2 _12710_ (.A(_07107_),
    .X(_07109_));
 sky130_fd_sc_hd__nor2_4 _12711_ (.A(\CPU_Xreg_value_a4[3][31] ),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__a211o_4 _12712_ (.A1(_06984_),
    .A2(_07108_),
    .B1(_07084_),
    .C1(_07110_),
    .X(_07111_));
 sky130_fd_sc_hd__inv_2 _12713_ (.A(_07111_),
    .Y(_00941_));
 sky130_fd_sc_hd__buf_2 _12714_ (.A(_07041_),
    .X(_07112_));
 sky130_fd_sc_hd__nor2_4 _12715_ (.A(\CPU_Xreg_value_a4[3][30] ),
    .B(_07109_),
    .Y(_07113_));
 sky130_fd_sc_hd__a211o_4 _12716_ (.A1(_06994_),
    .A2(_07108_),
    .B1(_07112_),
    .C1(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__inv_2 _12717_ (.A(_07114_),
    .Y(_00940_));
 sky130_fd_sc_hd__buf_2 _12718_ (.A(_07106_),
    .X(_07115_));
 sky130_fd_sc_hd__buf_2 _12719_ (.A(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__buf_2 _12720_ (.A(_07107_),
    .X(_07117_));
 sky130_fd_sc_hd__nor2_4 _12721_ (.A(\CPU_Xreg_value_a4[3][29] ),
    .B(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__a211o_4 _12722_ (.A1(_06997_),
    .A2(_07116_),
    .B1(_07112_),
    .C1(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__inv_2 _12723_ (.A(_07119_),
    .Y(_00939_));
 sky130_fd_sc_hd__nor2_4 _12724_ (.A(\CPU_Xreg_value_a4[3][28] ),
    .B(_07117_),
    .Y(_07120_));
 sky130_fd_sc_hd__a211o_4 _12725_ (.A1(_07001_),
    .A2(_07116_),
    .B1(_07112_),
    .C1(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__inv_2 _12726_ (.A(_07121_),
    .Y(_00938_));
 sky130_fd_sc_hd__nor2_4 _12727_ (.A(\CPU_Xreg_value_a4[3][27] ),
    .B(_07117_),
    .Y(_07122_));
 sky130_fd_sc_hd__a211o_4 _12728_ (.A1(_07005_),
    .A2(_07116_),
    .B1(_07112_),
    .C1(_07122_),
    .X(_07123_));
 sky130_fd_sc_hd__inv_2 _12729_ (.A(_07123_),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2_4 _12730_ (.A(\CPU_Xreg_value_a4[3][26] ),
    .B(_07117_),
    .Y(_07124_));
 sky130_fd_sc_hd__a211o_4 _12731_ (.A1(_07010_),
    .A2(_07116_),
    .B1(_07112_),
    .C1(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__inv_2 _12732_ (.A(_07125_),
    .Y(_00936_));
 sky130_fd_sc_hd__nor2_4 _12733_ (.A(\CPU_Xreg_value_a4[3][25] ),
    .B(_07117_),
    .Y(_07126_));
 sky130_fd_sc_hd__a211o_4 _12734_ (.A1(_07013_),
    .A2(_07116_),
    .B1(_07112_),
    .C1(_07126_),
    .X(_07127_));
 sky130_fd_sc_hd__inv_2 _12735_ (.A(_07127_),
    .Y(_00935_));
 sky130_fd_sc_hd__buf_2 _12736_ (.A(_07041_),
    .X(_07128_));
 sky130_fd_sc_hd__nor2_4 _12737_ (.A(\CPU_Xreg_value_a4[3][24] ),
    .B(_07117_),
    .Y(_07129_));
 sky130_fd_sc_hd__a211o_4 _12738_ (.A1(_07016_),
    .A2(_07116_),
    .B1(_07128_),
    .C1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__inv_2 _12739_ (.A(_07130_),
    .Y(_00934_));
 sky130_fd_sc_hd__buf_2 _12740_ (.A(_07115_),
    .X(_07131_));
 sky130_fd_sc_hd__buf_2 _12741_ (.A(_07107_),
    .X(_07132_));
 sky130_fd_sc_hd__nor2_4 _12742_ (.A(\CPU_Xreg_value_a4[3][23] ),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__a211o_4 _12743_ (.A1(_07019_),
    .A2(_07131_),
    .B1(_07128_),
    .C1(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__inv_2 _12744_ (.A(_07134_),
    .Y(_00933_));
 sky130_fd_sc_hd__nor2_4 _12745_ (.A(\CPU_Xreg_value_a4[3][22] ),
    .B(_07132_),
    .Y(_07135_));
 sky130_fd_sc_hd__a211o_4 _12746_ (.A1(_07023_),
    .A2(_07131_),
    .B1(_07128_),
    .C1(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__inv_2 _12747_ (.A(_07136_),
    .Y(_00932_));
 sky130_fd_sc_hd__nor2_4 _12748_ (.A(\CPU_Xreg_value_a4[3][21] ),
    .B(_07132_),
    .Y(_07137_));
 sky130_fd_sc_hd__a211o_4 _12749_ (.A1(_07027_),
    .A2(_07131_),
    .B1(_07128_),
    .C1(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__inv_2 _12750_ (.A(_07138_),
    .Y(_00931_));
 sky130_fd_sc_hd__nor2_4 _12751_ (.A(\CPU_Xreg_value_a4[3][20] ),
    .B(_07132_),
    .Y(_07139_));
 sky130_fd_sc_hd__a211o_4 _12752_ (.A1(_07031_),
    .A2(_07131_),
    .B1(_07128_),
    .C1(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__inv_2 _12753_ (.A(_07140_),
    .Y(_00930_));
 sky130_fd_sc_hd__nor2_4 _12754_ (.A(\CPU_Xreg_value_a4[3][19] ),
    .B(_07132_),
    .Y(_07141_));
 sky130_fd_sc_hd__a211o_4 _12755_ (.A1(_07034_),
    .A2(_07131_),
    .B1(_07128_),
    .C1(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__inv_2 _12756_ (.A(_07142_),
    .Y(_00929_));
 sky130_fd_sc_hd__buf_2 _12757_ (.A(_07041_),
    .X(_07143_));
 sky130_fd_sc_hd__nor2_4 _12758_ (.A(\CPU_Xreg_value_a4[3][18] ),
    .B(_07132_),
    .Y(_07144_));
 sky130_fd_sc_hd__a211o_4 _12759_ (.A1(_07037_),
    .A2(_07131_),
    .B1(_07143_),
    .C1(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__inv_2 _12760_ (.A(_07145_),
    .Y(_00928_));
 sky130_fd_sc_hd__buf_2 _12761_ (.A(_07107_),
    .X(_07146_));
 sky130_fd_sc_hd__buf_2 _12762_ (.A(_07106_),
    .X(_07147_));
 sky130_fd_sc_hd__nor2_4 _12763_ (.A(\CPU_Xreg_value_a4[3][17] ),
    .B(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__a211o_4 _12764_ (.A1(_07040_),
    .A2(_07146_),
    .B1(_07143_),
    .C1(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__inv_2 _12765_ (.A(_07149_),
    .Y(_00927_));
 sky130_fd_sc_hd__nor2_4 _12766_ (.A(\CPU_Xreg_value_a4[3][16] ),
    .B(_07147_),
    .Y(_07150_));
 sky130_fd_sc_hd__a211o_4 _12767_ (.A1(_07045_),
    .A2(_07146_),
    .B1(_07143_),
    .C1(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__inv_2 _12768_ (.A(_07151_),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_4 _12769_ (.A(\CPU_Xreg_value_a4[3][15] ),
    .B(_07147_),
    .Y(_07152_));
 sky130_fd_sc_hd__a211o_4 _12770_ (.A1(_07049_),
    .A2(_07146_),
    .B1(_07143_),
    .C1(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__inv_2 _12771_ (.A(_07153_),
    .Y(_00925_));
 sky130_fd_sc_hd__nor2_4 _12772_ (.A(\CPU_Xreg_value_a4[3][14] ),
    .B(_07147_),
    .Y(_07154_));
 sky130_fd_sc_hd__a211o_4 _12773_ (.A1(_07053_),
    .A2(_07146_),
    .B1(_07143_),
    .C1(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__inv_2 _12774_ (.A(_07155_),
    .Y(_00924_));
 sky130_fd_sc_hd__nor2_4 _12775_ (.A(\CPU_Xreg_value_a4[3][13] ),
    .B(_07147_),
    .Y(_07156_));
 sky130_fd_sc_hd__a211o_4 _12776_ (.A1(_07056_),
    .A2(_07146_),
    .B1(_07143_),
    .C1(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__inv_2 _12777_ (.A(_07157_),
    .Y(_00923_));
 sky130_fd_sc_hd__buf_2 _12778_ (.A(CPU_reset_a3),
    .X(_07158_));
 sky130_fd_sc_hd__buf_2 _12779_ (.A(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__buf_2 _12780_ (.A(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__nor2_4 _12781_ (.A(\CPU_Xreg_value_a4[3][12] ),
    .B(_07147_),
    .Y(_07161_));
 sky130_fd_sc_hd__a211o_4 _12782_ (.A1(_07059_),
    .A2(_07146_),
    .B1(_07160_),
    .C1(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__inv_2 _12783_ (.A(_07162_),
    .Y(_00922_));
 sky130_fd_sc_hd__buf_2 _12784_ (.A(_07107_),
    .X(_07163_));
 sky130_fd_sc_hd__buf_2 _12785_ (.A(_07106_),
    .X(_07164_));
 sky130_fd_sc_hd__nor2_4 _12786_ (.A(\CPU_Xreg_value_a4[3][11] ),
    .B(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__a211o_4 _12787_ (.A1(_07062_),
    .A2(_07163_),
    .B1(_07160_),
    .C1(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__inv_2 _12788_ (.A(_07166_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_4 _12789_ (.A(\CPU_Xreg_value_a4[3][10] ),
    .B(_07164_),
    .Y(_07167_));
 sky130_fd_sc_hd__a211o_4 _12790_ (.A1(_07066_),
    .A2(_07163_),
    .B1(_07160_),
    .C1(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__inv_2 _12791_ (.A(_07168_),
    .Y(_00920_));
 sky130_fd_sc_hd__nor2_4 _12792_ (.A(\CPU_Xreg_value_a4[3][9] ),
    .B(_07164_),
    .Y(_07169_));
 sky130_fd_sc_hd__a211o_4 _12793_ (.A1(_07070_),
    .A2(_07163_),
    .B1(_07160_),
    .C1(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__inv_2 _12794_ (.A(_07170_),
    .Y(_00919_));
 sky130_fd_sc_hd__nor2_4 _12795_ (.A(\CPU_Xreg_value_a4[3][8] ),
    .B(_07164_),
    .Y(_07171_));
 sky130_fd_sc_hd__a211o_4 _12796_ (.A1(_07074_),
    .A2(_07163_),
    .B1(_07160_),
    .C1(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__inv_2 _12797_ (.A(_07172_),
    .Y(_00918_));
 sky130_fd_sc_hd__nor2_4 _12798_ (.A(\CPU_Xreg_value_a4[3][7] ),
    .B(_07164_),
    .Y(_07173_));
 sky130_fd_sc_hd__a211o_4 _12799_ (.A1(_07077_),
    .A2(_07163_),
    .B1(_07160_),
    .C1(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__inv_2 _12800_ (.A(_07174_),
    .Y(_00917_));
 sky130_fd_sc_hd__buf_2 _12801_ (.A(_07159_),
    .X(_07175_));
 sky130_fd_sc_hd__nor2_4 _12802_ (.A(\CPU_Xreg_value_a4[3][6] ),
    .B(_07164_),
    .Y(_07176_));
 sky130_fd_sc_hd__a211o_4 _12803_ (.A1(_07080_),
    .A2(_07163_),
    .B1(_07175_),
    .C1(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__inv_2 _12804_ (.A(_07177_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_4 _12805_ (.A(\CPU_Xreg_value_a4[3][5] ),
    .B(_07115_),
    .Y(_07178_));
 sky130_fd_sc_hd__a211o_4 _12806_ (.A1(_07083_),
    .A2(_07109_),
    .B1(_07175_),
    .C1(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__inv_2 _12807_ (.A(_07179_),
    .Y(_00915_));
 sky130_fd_sc_hd__nor2_4 _12808_ (.A(\CPU_Xreg_value_a4[3][4] ),
    .B(_07115_),
    .Y(_07180_));
 sky130_fd_sc_hd__a211o_4 _12809_ (.A1(_07087_),
    .A2(_07109_),
    .B1(_07175_),
    .C1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__inv_2 _12810_ (.A(_07181_),
    .Y(_00914_));
 sky130_fd_sc_hd__nor2_4 _12811_ (.A(\CPU_Xreg_value_a4[3][3] ),
    .B(_07115_),
    .Y(_07182_));
 sky130_fd_sc_hd__a211o_4 _12812_ (.A1(_07090_),
    .A2(_07109_),
    .B1(_07175_),
    .C1(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__inv_2 _12813_ (.A(_07183_),
    .Y(_00913_));
 sky130_fd_sc_hd__nor2_4 _12814_ (.A(\CPU_Xreg_value_a4[3][2] ),
    .B(_07115_),
    .Y(_07184_));
 sky130_fd_sc_hd__a211o_4 _12815_ (.A1(_07093_),
    .A2(_07109_),
    .B1(_07175_),
    .C1(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__inv_2 _12816_ (.A(_07185_),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _12817_ (.A(\CPU_Xreg_value_a4[3][1] ),
    .Y(_07186_));
 sky130_fd_sc_hd__nor2_4 _12818_ (.A(_07186_),
    .B(_07108_),
    .Y(_07187_));
 sky130_fd_sc_hd__a211o_4 _12819_ (.A1(_07097_),
    .A2(_07108_),
    .B1(_06140_),
    .C1(_07187_),
    .X(_00911_));
 sky130_fd_sc_hd__buf_2 _12820_ (.A(_06981_),
    .X(_07188_));
 sky130_fd_sc_hd__inv_2 _12821_ (.A(\CPU_Xreg_value_a4[3][0] ),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_4 _12822_ (.A(_07189_),
    .B(_07108_),
    .Y(_07190_));
 sky130_fd_sc_hd__a211o_4 _12823_ (.A1(_07188_),
    .A2(_07108_),
    .B1(_06140_),
    .C1(_07190_),
    .X(_00910_));
 sky130_fd_sc_hd__inv_2 _12824_ (.A(_06145_),
    .Y(_07191_));
 sky130_fd_sc_hd__or2_4 _12825_ (.A(_07191_),
    .B(_06147_),
    .X(_07192_));
 sky130_fd_sc_hd__or2_4 _12826_ (.A(_06156_),
    .B(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__nor2_4 _12827_ (.A(_06166_),
    .B(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__buf_2 _12828_ (.A(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__buf_2 _12829_ (.A(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__buf_2 _12830_ (.A(_07195_),
    .X(_07197_));
 sky130_fd_sc_hd__nor2_4 _12831_ (.A(\CPU_Xreg_value_a4[4][31] ),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__a211o_4 _12832_ (.A1(_06984_),
    .A2(_07196_),
    .B1(_07175_),
    .C1(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__inv_2 _12833_ (.A(_07199_),
    .Y(_00909_));
 sky130_fd_sc_hd__buf_2 _12834_ (.A(_07159_),
    .X(_07200_));
 sky130_fd_sc_hd__nor2_4 _12835_ (.A(\CPU_Xreg_value_a4[4][30] ),
    .B(_07197_),
    .Y(_07201_));
 sky130_fd_sc_hd__a211o_4 _12836_ (.A1(_06994_),
    .A2(_07196_),
    .B1(_07200_),
    .C1(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__inv_2 _12837_ (.A(_07202_),
    .Y(_00908_));
 sky130_fd_sc_hd__nor2_4 _12838_ (.A(\CPU_Xreg_value_a4[4][29] ),
    .B(_07197_),
    .Y(_07203_));
 sky130_fd_sc_hd__a211o_4 _12839_ (.A1(_06997_),
    .A2(_07196_),
    .B1(_07200_),
    .C1(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__inv_2 _12840_ (.A(_07204_),
    .Y(_00907_));
 sky130_fd_sc_hd__buf_2 _12841_ (.A(_07195_),
    .X(_07205_));
 sky130_fd_sc_hd__nor2_4 _12842_ (.A(\CPU_Xreg_value_a4[4][28] ),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__a211o_4 _12843_ (.A1(_07001_),
    .A2(_07196_),
    .B1(_07200_),
    .C1(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__inv_2 _12844_ (.A(_07207_),
    .Y(_00906_));
 sky130_fd_sc_hd__buf_2 _12845_ (.A(_07194_),
    .X(_07208_));
 sky130_fd_sc_hd__buf_2 _12846_ (.A(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__nor2_4 _12847_ (.A(\CPU_Xreg_value_a4[4][27] ),
    .B(_07205_),
    .Y(_07210_));
 sky130_fd_sc_hd__a211o_4 _12848_ (.A1(_07005_),
    .A2(_07209_),
    .B1(_07200_),
    .C1(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__inv_2 _12849_ (.A(_07211_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_4 _12850_ (.A(\CPU_Xreg_value_a4[4][26] ),
    .B(_07205_),
    .Y(_07212_));
 sky130_fd_sc_hd__a211o_4 _12851_ (.A1(_07010_),
    .A2(_07209_),
    .B1(_07200_),
    .C1(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__inv_2 _12852_ (.A(_07213_),
    .Y(_00904_));
 sky130_fd_sc_hd__nor2_4 _12853_ (.A(\CPU_Xreg_value_a4[4][25] ),
    .B(_07205_),
    .Y(_07214_));
 sky130_fd_sc_hd__a211o_4 _12854_ (.A1(_07013_),
    .A2(_07209_),
    .B1(_07200_),
    .C1(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__inv_2 _12855_ (.A(_07215_),
    .Y(_00903_));
 sky130_fd_sc_hd__buf_2 _12856_ (.A(_07159_),
    .X(_07216_));
 sky130_fd_sc_hd__nor2_4 _12857_ (.A(\CPU_Xreg_value_a4[4][24] ),
    .B(_07205_),
    .Y(_07217_));
 sky130_fd_sc_hd__a211o_4 _12858_ (.A1(_07016_),
    .A2(_07209_),
    .B1(_07216_),
    .C1(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__inv_2 _12859_ (.A(_07218_),
    .Y(_00902_));
 sky130_fd_sc_hd__nor2_4 _12860_ (.A(\CPU_Xreg_value_a4[4][23] ),
    .B(_07205_),
    .Y(_07219_));
 sky130_fd_sc_hd__a211o_4 _12861_ (.A1(_07019_),
    .A2(_07209_),
    .B1(_07216_),
    .C1(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__inv_2 _12862_ (.A(_07220_),
    .Y(_00901_));
 sky130_fd_sc_hd__buf_2 _12863_ (.A(_07195_),
    .X(_07221_));
 sky130_fd_sc_hd__nor2_4 _12864_ (.A(\CPU_Xreg_value_a4[4][22] ),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__a211o_4 _12865_ (.A1(_07023_),
    .A2(_07209_),
    .B1(_07216_),
    .C1(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__inv_2 _12866_ (.A(_07223_),
    .Y(_00900_));
 sky130_fd_sc_hd__buf_2 _12867_ (.A(_07208_),
    .X(_07224_));
 sky130_fd_sc_hd__nor2_4 _12868_ (.A(\CPU_Xreg_value_a4[4][21] ),
    .B(_07221_),
    .Y(_07225_));
 sky130_fd_sc_hd__a211o_4 _12869_ (.A1(_07027_),
    .A2(_07224_),
    .B1(_07216_),
    .C1(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__inv_2 _12870_ (.A(_07226_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_4 _12871_ (.A(\CPU_Xreg_value_a4[4][20] ),
    .B(_07221_),
    .Y(_07227_));
 sky130_fd_sc_hd__a211o_4 _12872_ (.A1(_07031_),
    .A2(_07224_),
    .B1(_07216_),
    .C1(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__inv_2 _12873_ (.A(_07228_),
    .Y(_00898_));
 sky130_fd_sc_hd__nor2_4 _12874_ (.A(\CPU_Xreg_value_a4[4][19] ),
    .B(_07221_),
    .Y(_07229_));
 sky130_fd_sc_hd__a211o_4 _12875_ (.A1(_07034_),
    .A2(_07224_),
    .B1(_07216_),
    .C1(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__inv_2 _12876_ (.A(_07230_),
    .Y(_00897_));
 sky130_fd_sc_hd__buf_2 _12877_ (.A(_07159_),
    .X(_07231_));
 sky130_fd_sc_hd__nor2_4 _12878_ (.A(\CPU_Xreg_value_a4[4][18] ),
    .B(_07221_),
    .Y(_07232_));
 sky130_fd_sc_hd__a211o_4 _12879_ (.A1(_07037_),
    .A2(_07224_),
    .B1(_07231_),
    .C1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__inv_2 _12880_ (.A(_07233_),
    .Y(_00896_));
 sky130_fd_sc_hd__nor2_4 _12881_ (.A(\CPU_Xreg_value_a4[4][17] ),
    .B(_07221_),
    .Y(_07234_));
 sky130_fd_sc_hd__a211o_4 _12882_ (.A1(_07040_),
    .A2(_07224_),
    .B1(_07231_),
    .C1(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__inv_2 _12883_ (.A(_07235_),
    .Y(_00895_));
 sky130_fd_sc_hd__buf_2 _12884_ (.A(_07194_),
    .X(_07236_));
 sky130_fd_sc_hd__nor2_4 _12885_ (.A(\CPU_Xreg_value_a4[4][16] ),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__a211o_4 _12886_ (.A1(_07045_),
    .A2(_07224_),
    .B1(_07231_),
    .C1(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__inv_2 _12887_ (.A(_07238_),
    .Y(_00894_));
 sky130_fd_sc_hd__buf_2 _12888_ (.A(_07195_),
    .X(_07239_));
 sky130_fd_sc_hd__nor2_4 _12889_ (.A(\CPU_Xreg_value_a4[4][15] ),
    .B(_07236_),
    .Y(_07240_));
 sky130_fd_sc_hd__a211o_4 _12890_ (.A1(_07049_),
    .A2(_07239_),
    .B1(_07231_),
    .C1(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(_07241_),
    .Y(_00893_));
 sky130_fd_sc_hd__nor2_4 _12892_ (.A(\CPU_Xreg_value_a4[4][14] ),
    .B(_07236_),
    .Y(_07242_));
 sky130_fd_sc_hd__a211o_4 _12893_ (.A1(_07053_),
    .A2(_07239_),
    .B1(_07231_),
    .C1(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__inv_2 _12894_ (.A(_07243_),
    .Y(_00892_));
 sky130_fd_sc_hd__nor2_4 _12895_ (.A(\CPU_Xreg_value_a4[4][13] ),
    .B(_07236_),
    .Y(_07244_));
 sky130_fd_sc_hd__a211o_4 _12896_ (.A1(_07056_),
    .A2(_07239_),
    .B1(_07231_),
    .C1(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__inv_2 _12897_ (.A(_07245_),
    .Y(_00891_));
 sky130_fd_sc_hd__buf_2 _12898_ (.A(_07159_),
    .X(_07246_));
 sky130_fd_sc_hd__nor2_4 _12899_ (.A(\CPU_Xreg_value_a4[4][12] ),
    .B(_07236_),
    .Y(_07247_));
 sky130_fd_sc_hd__a211o_4 _12900_ (.A1(_07059_),
    .A2(_07239_),
    .B1(_07246_),
    .C1(_07247_),
    .X(_07248_));
 sky130_fd_sc_hd__inv_2 _12901_ (.A(_07248_),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_4 _12902_ (.A(\CPU_Xreg_value_a4[4][11] ),
    .B(_07236_),
    .Y(_07249_));
 sky130_fd_sc_hd__a211o_4 _12903_ (.A1(_07062_),
    .A2(_07239_),
    .B1(_07246_),
    .C1(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__inv_2 _12904_ (.A(_07250_),
    .Y(_00889_));
 sky130_fd_sc_hd__buf_2 _12905_ (.A(_07194_),
    .X(_07251_));
 sky130_fd_sc_hd__nor2_4 _12906_ (.A(\CPU_Xreg_value_a4[4][10] ),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__a211o_4 _12907_ (.A1(_07066_),
    .A2(_07239_),
    .B1(_07246_),
    .C1(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__inv_2 _12908_ (.A(_07253_),
    .Y(_00888_));
 sky130_fd_sc_hd__buf_2 _12909_ (.A(_07195_),
    .X(_07254_));
 sky130_fd_sc_hd__nor2_4 _12910_ (.A(\CPU_Xreg_value_a4[4][9] ),
    .B(_07251_),
    .Y(_07255_));
 sky130_fd_sc_hd__a211o_4 _12911_ (.A1(_07070_),
    .A2(_07254_),
    .B1(_07246_),
    .C1(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__inv_2 _12912_ (.A(_07256_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_4 _12913_ (.A(\CPU_Xreg_value_a4[4][8] ),
    .B(_07251_),
    .Y(_07257_));
 sky130_fd_sc_hd__a211o_4 _12914_ (.A1(_07074_),
    .A2(_07254_),
    .B1(_07246_),
    .C1(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__inv_2 _12915_ (.A(_07258_),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_4 _12916_ (.A(\CPU_Xreg_value_a4[4][7] ),
    .B(_07251_),
    .Y(_07259_));
 sky130_fd_sc_hd__a211o_4 _12917_ (.A1(_07077_),
    .A2(_07254_),
    .B1(_07246_),
    .C1(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__inv_2 _12918_ (.A(_07260_),
    .Y(_00885_));
 sky130_fd_sc_hd__buf_2 _12919_ (.A(_07158_),
    .X(_07261_));
 sky130_fd_sc_hd__buf_2 _12920_ (.A(_07261_),
    .X(_07262_));
 sky130_fd_sc_hd__nor2_4 _12921_ (.A(\CPU_Xreg_value_a4[4][6] ),
    .B(_07251_),
    .Y(_07263_));
 sky130_fd_sc_hd__a211o_4 _12922_ (.A1(_07080_),
    .A2(_07254_),
    .B1(_07262_),
    .C1(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__inv_2 _12923_ (.A(_07264_),
    .Y(_00884_));
 sky130_fd_sc_hd__nor2_4 _12924_ (.A(\CPU_Xreg_value_a4[4][5] ),
    .B(_07251_),
    .Y(_07265_));
 sky130_fd_sc_hd__a211o_4 _12925_ (.A1(_07083_),
    .A2(_07254_),
    .B1(_07262_),
    .C1(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__inv_2 _12926_ (.A(_07266_),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2_4 _12927_ (.A(\CPU_Xreg_value_a4[4][4] ),
    .B(_07208_),
    .Y(_07267_));
 sky130_fd_sc_hd__a211o_4 _12928_ (.A1(_07087_),
    .A2(_07254_),
    .B1(_07262_),
    .C1(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__inv_2 _12929_ (.A(_07268_),
    .Y(_00882_));
 sky130_fd_sc_hd__nor2_4 _12930_ (.A(\CPU_Xreg_value_a4[4][3] ),
    .B(_07208_),
    .Y(_07269_));
 sky130_fd_sc_hd__a211o_4 _12931_ (.A1(_07090_),
    .A2(_07197_),
    .B1(_07262_),
    .C1(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(_07270_),
    .Y(_00881_));
 sky130_fd_sc_hd__buf_2 _12933_ (.A(_06859_),
    .X(_07271_));
 sky130_fd_sc_hd__buf_2 _12934_ (.A(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__buf_2 _12935_ (.A(_06101_),
    .X(_07273_));
 sky130_fd_sc_hd__buf_2 _12936_ (.A(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__inv_2 _12937_ (.A(\CPU_Xreg_value_a4[4][2] ),
    .Y(_07275_));
 sky130_fd_sc_hd__nor2_4 _12938_ (.A(_07275_),
    .B(_07196_),
    .Y(_07276_));
 sky130_fd_sc_hd__a211o_4 _12939_ (.A1(_07272_),
    .A2(_07196_),
    .B1(_07274_),
    .C1(_07276_),
    .X(_00880_));
 sky130_fd_sc_hd__buf_2 _12940_ (.A(_06868_),
    .X(_07277_));
 sky130_fd_sc_hd__nor2_4 _12941_ (.A(\CPU_Xreg_value_a4[4][1] ),
    .B(_07208_),
    .Y(_07278_));
 sky130_fd_sc_hd__a211o_4 _12942_ (.A1(_07277_),
    .A2(_07197_),
    .B1(_07262_),
    .C1(_07278_),
    .X(_07279_));
 sky130_fd_sc_hd__inv_2 _12943_ (.A(_07279_),
    .Y(_00879_));
 sky130_fd_sc_hd__nor2_4 _12944_ (.A(\CPU_Xreg_value_a4[4][0] ),
    .B(_07208_),
    .Y(_07280_));
 sky130_fd_sc_hd__a211o_4 _12945_ (.A1(_07101_),
    .A2(_07197_),
    .B1(_07262_),
    .C1(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__inv_2 _12946_ (.A(_07281_),
    .Y(_00878_));
 sky130_fd_sc_hd__or2_4 _12947_ (.A(_06152_),
    .B(_07192_),
    .X(_07282_));
 sky130_fd_sc_hd__nor2_4 _12948_ (.A(_06166_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__buf_2 _12949_ (.A(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__buf_2 _12950_ (.A(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__buf_2 _12951_ (.A(_07261_),
    .X(_07286_));
 sky130_fd_sc_hd__buf_2 _12952_ (.A(_07284_),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_4 _12953_ (.A(\CPU_Xreg_value_a4[5][31] ),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__a211o_4 _12954_ (.A1(_06984_),
    .A2(_07285_),
    .B1(_07286_),
    .C1(_07288_),
    .X(_07289_));
 sky130_fd_sc_hd__inv_2 _12955_ (.A(_07289_),
    .Y(_00877_));
 sky130_fd_sc_hd__nor2_4 _12956_ (.A(\CPU_Xreg_value_a4[5][30] ),
    .B(_07287_),
    .Y(_07290_));
 sky130_fd_sc_hd__a211o_4 _12957_ (.A1(_06994_),
    .A2(_07285_),
    .B1(_07286_),
    .C1(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__inv_2 _12958_ (.A(_07291_),
    .Y(_00876_));
 sky130_fd_sc_hd__buf_2 _12959_ (.A(_07283_),
    .X(_07292_));
 sky130_fd_sc_hd__buf_2 _12960_ (.A(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__buf_2 _12961_ (.A(_07284_),
    .X(_07294_));
 sky130_fd_sc_hd__nor2_4 _12962_ (.A(\CPU_Xreg_value_a4[5][29] ),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__a211o_4 _12963_ (.A1(_06997_),
    .A2(_07293_),
    .B1(_07286_),
    .C1(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__inv_2 _12964_ (.A(_07296_),
    .Y(_00875_));
 sky130_fd_sc_hd__nor2_4 _12965_ (.A(\CPU_Xreg_value_a4[5][28] ),
    .B(_07294_),
    .Y(_07297_));
 sky130_fd_sc_hd__a211o_4 _12966_ (.A1(_07001_),
    .A2(_07293_),
    .B1(_07286_),
    .C1(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__inv_2 _12967_ (.A(_07298_),
    .Y(_00874_));
 sky130_fd_sc_hd__nor2_4 _12968_ (.A(\CPU_Xreg_value_a4[5][27] ),
    .B(_07294_),
    .Y(_07299_));
 sky130_fd_sc_hd__a211o_4 _12969_ (.A1(_07005_),
    .A2(_07293_),
    .B1(_07286_),
    .C1(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__inv_2 _12970_ (.A(_07300_),
    .Y(_00873_));
 sky130_fd_sc_hd__nor2_4 _12971_ (.A(\CPU_Xreg_value_a4[5][26] ),
    .B(_07294_),
    .Y(_07301_));
 sky130_fd_sc_hd__a211o_4 _12972_ (.A1(_07010_),
    .A2(_07293_),
    .B1(_07286_),
    .C1(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__inv_2 _12973_ (.A(_07302_),
    .Y(_00872_));
 sky130_fd_sc_hd__buf_2 _12974_ (.A(_07261_),
    .X(_07303_));
 sky130_fd_sc_hd__nor2_4 _12975_ (.A(\CPU_Xreg_value_a4[5][25] ),
    .B(_07294_),
    .Y(_07304_));
 sky130_fd_sc_hd__a211o_4 _12976_ (.A1(_07013_),
    .A2(_07293_),
    .B1(_07303_),
    .C1(_07304_),
    .X(_07305_));
 sky130_fd_sc_hd__inv_2 _12977_ (.A(_07305_),
    .Y(_00871_));
 sky130_fd_sc_hd__nor2_4 _12978_ (.A(\CPU_Xreg_value_a4[5][24] ),
    .B(_07294_),
    .Y(_07306_));
 sky130_fd_sc_hd__a211o_4 _12979_ (.A1(_07016_),
    .A2(_07293_),
    .B1(_07303_),
    .C1(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__inv_2 _12980_ (.A(_07307_),
    .Y(_00870_));
 sky130_fd_sc_hd__buf_2 _12981_ (.A(_07292_),
    .X(_07308_));
 sky130_fd_sc_hd__buf_2 _12982_ (.A(_07284_),
    .X(_07309_));
 sky130_fd_sc_hd__nor2_4 _12983_ (.A(\CPU_Xreg_value_a4[5][23] ),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__a211o_4 _12984_ (.A1(_07019_),
    .A2(_07308_),
    .B1(_07303_),
    .C1(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__inv_2 _12985_ (.A(_07311_),
    .Y(_00869_));
 sky130_fd_sc_hd__nor2_4 _12986_ (.A(\CPU_Xreg_value_a4[5][22] ),
    .B(_07309_),
    .Y(_07312_));
 sky130_fd_sc_hd__a211o_4 _12987_ (.A1(_07023_),
    .A2(_07308_),
    .B1(_07303_),
    .C1(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__inv_2 _12988_ (.A(_07313_),
    .Y(_00868_));
 sky130_fd_sc_hd__nor2_4 _12989_ (.A(\CPU_Xreg_value_a4[5][21] ),
    .B(_07309_),
    .Y(_07314_));
 sky130_fd_sc_hd__a211o_4 _12990_ (.A1(_07027_),
    .A2(_07308_),
    .B1(_07303_),
    .C1(_07314_),
    .X(_07315_));
 sky130_fd_sc_hd__inv_2 _12991_ (.A(_07315_),
    .Y(_00867_));
 sky130_fd_sc_hd__nor2_4 _12992_ (.A(\CPU_Xreg_value_a4[5][20] ),
    .B(_07309_),
    .Y(_07316_));
 sky130_fd_sc_hd__a211o_4 _12993_ (.A1(_07031_),
    .A2(_07308_),
    .B1(_07303_),
    .C1(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__inv_2 _12994_ (.A(_07317_),
    .Y(_00866_));
 sky130_fd_sc_hd__buf_2 _12995_ (.A(_07261_),
    .X(_07318_));
 sky130_fd_sc_hd__nor2_4 _12996_ (.A(\CPU_Xreg_value_a4[5][19] ),
    .B(_07309_),
    .Y(_07319_));
 sky130_fd_sc_hd__a211o_4 _12997_ (.A1(_07034_),
    .A2(_07308_),
    .B1(_07318_),
    .C1(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__inv_2 _12998_ (.A(_07320_),
    .Y(_00865_));
 sky130_fd_sc_hd__nor2_4 _12999_ (.A(\CPU_Xreg_value_a4[5][18] ),
    .B(_07309_),
    .Y(_07321_));
 sky130_fd_sc_hd__a211o_4 _13000_ (.A1(_07037_),
    .A2(_07308_),
    .B1(_07318_),
    .C1(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__inv_2 _13001_ (.A(_07322_),
    .Y(_00864_));
 sky130_fd_sc_hd__buf_2 _13002_ (.A(_07284_),
    .X(_07323_));
 sky130_fd_sc_hd__buf_2 _13003_ (.A(_07283_),
    .X(_07324_));
 sky130_fd_sc_hd__nor2_4 _13004_ (.A(\CPU_Xreg_value_a4[5][17] ),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__a211o_4 _13005_ (.A1(_07040_),
    .A2(_07323_),
    .B1(_07318_),
    .C1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__inv_2 _13006_ (.A(_07326_),
    .Y(_00863_));
 sky130_fd_sc_hd__nor2_4 _13007_ (.A(\CPU_Xreg_value_a4[5][16] ),
    .B(_07324_),
    .Y(_07327_));
 sky130_fd_sc_hd__a211o_4 _13008_ (.A1(_07045_),
    .A2(_07323_),
    .B1(_07318_),
    .C1(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__inv_2 _13009_ (.A(_07328_),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_4 _13010_ (.A(\CPU_Xreg_value_a4[5][15] ),
    .B(_07324_),
    .Y(_07329_));
 sky130_fd_sc_hd__a211o_4 _13011_ (.A1(_07049_),
    .A2(_07323_),
    .B1(_07318_),
    .C1(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__inv_2 _13012_ (.A(_07330_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor2_4 _13013_ (.A(\CPU_Xreg_value_a4[5][14] ),
    .B(_07324_),
    .Y(_07331_));
 sky130_fd_sc_hd__a211o_4 _13014_ (.A1(_07053_),
    .A2(_07323_),
    .B1(_07318_),
    .C1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__inv_2 _13015_ (.A(_07332_),
    .Y(_00860_));
 sky130_fd_sc_hd__buf_2 _13016_ (.A(_07261_),
    .X(_07333_));
 sky130_fd_sc_hd__nor2_4 _13017_ (.A(\CPU_Xreg_value_a4[5][13] ),
    .B(_07324_),
    .Y(_07334_));
 sky130_fd_sc_hd__a211o_4 _13018_ (.A1(_07056_),
    .A2(_07323_),
    .B1(_07333_),
    .C1(_07334_),
    .X(_07335_));
 sky130_fd_sc_hd__inv_2 _13019_ (.A(_07335_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor2_4 _13020_ (.A(\CPU_Xreg_value_a4[5][12] ),
    .B(_07324_),
    .Y(_07336_));
 sky130_fd_sc_hd__a211o_4 _13021_ (.A1(_07059_),
    .A2(_07323_),
    .B1(_07333_),
    .C1(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__inv_2 _13022_ (.A(_07337_),
    .Y(_00858_));
 sky130_fd_sc_hd__buf_2 _13023_ (.A(_07284_),
    .X(_07338_));
 sky130_fd_sc_hd__buf_2 _13024_ (.A(_07283_),
    .X(_07339_));
 sky130_fd_sc_hd__nor2_4 _13025_ (.A(\CPU_Xreg_value_a4[5][11] ),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__a211o_4 _13026_ (.A1(_07062_),
    .A2(_07338_),
    .B1(_07333_),
    .C1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__inv_2 _13027_ (.A(_07341_),
    .Y(_00857_));
 sky130_fd_sc_hd__nor2_4 _13028_ (.A(\CPU_Xreg_value_a4[5][10] ),
    .B(_07339_),
    .Y(_07342_));
 sky130_fd_sc_hd__a211o_4 _13029_ (.A1(_07066_),
    .A2(_07338_),
    .B1(_07333_),
    .C1(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__inv_2 _13030_ (.A(_07343_),
    .Y(_00856_));
 sky130_fd_sc_hd__nor2_4 _13031_ (.A(\CPU_Xreg_value_a4[5][9] ),
    .B(_07339_),
    .Y(_07344_));
 sky130_fd_sc_hd__a211o_4 _13032_ (.A1(_07070_),
    .A2(_07338_),
    .B1(_07333_),
    .C1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__inv_2 _13033_ (.A(_07345_),
    .Y(_00855_));
 sky130_fd_sc_hd__nor2_4 _13034_ (.A(\CPU_Xreg_value_a4[5][8] ),
    .B(_07339_),
    .Y(_07346_));
 sky130_fd_sc_hd__a211o_4 _13035_ (.A1(_07074_),
    .A2(_07338_),
    .B1(_07333_),
    .C1(_07346_),
    .X(_07347_));
 sky130_fd_sc_hd__inv_2 _13036_ (.A(_07347_),
    .Y(_00854_));
 sky130_fd_sc_hd__buf_2 _13037_ (.A(_07261_),
    .X(_07348_));
 sky130_fd_sc_hd__nor2_4 _13038_ (.A(\CPU_Xreg_value_a4[5][7] ),
    .B(_07339_),
    .Y(_07349_));
 sky130_fd_sc_hd__a211o_4 _13039_ (.A1(_07077_),
    .A2(_07338_),
    .B1(_07348_),
    .C1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__inv_2 _13040_ (.A(_07350_),
    .Y(_00853_));
 sky130_fd_sc_hd__nor2_4 _13041_ (.A(\CPU_Xreg_value_a4[5][6] ),
    .B(_07339_),
    .Y(_07351_));
 sky130_fd_sc_hd__a211o_4 _13042_ (.A1(_07080_),
    .A2(_07338_),
    .B1(_07348_),
    .C1(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__inv_2 _13043_ (.A(_07352_),
    .Y(_00852_));
 sky130_fd_sc_hd__nor2_4 _13044_ (.A(\CPU_Xreg_value_a4[5][5] ),
    .B(_07292_),
    .Y(_07353_));
 sky130_fd_sc_hd__a211o_4 _13045_ (.A1(_07083_),
    .A2(_07287_),
    .B1(_07348_),
    .C1(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__inv_2 _13046_ (.A(_07354_),
    .Y(_00851_));
 sky130_fd_sc_hd__nor2_4 _13047_ (.A(\CPU_Xreg_value_a4[5][4] ),
    .B(_07292_),
    .Y(_07355_));
 sky130_fd_sc_hd__a211o_4 _13048_ (.A1(_07087_),
    .A2(_07287_),
    .B1(_07348_),
    .C1(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__inv_2 _13049_ (.A(_07356_),
    .Y(_00850_));
 sky130_fd_sc_hd__nor2_4 _13050_ (.A(\CPU_Xreg_value_a4[5][3] ),
    .B(_07292_),
    .Y(_07357_));
 sky130_fd_sc_hd__a211o_4 _13051_ (.A1(_07090_),
    .A2(_07287_),
    .B1(_07348_),
    .C1(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__inv_2 _13052_ (.A(_07358_),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _13053_ (.A(\CPU_Xreg_value_a4[5][2] ),
    .Y(_07359_));
 sky130_fd_sc_hd__nor2_4 _13054_ (.A(_07359_),
    .B(_07285_),
    .Y(_07360_));
 sky130_fd_sc_hd__a211o_4 _13055_ (.A1(_07272_),
    .A2(_07285_),
    .B1(_07274_),
    .C1(_07360_),
    .X(_00848_));
 sky130_fd_sc_hd__nor2_4 _13056_ (.A(\CPU_Xreg_value_a4[5][1] ),
    .B(_07292_),
    .Y(_07361_));
 sky130_fd_sc_hd__a211o_4 _13057_ (.A1(_07277_),
    .A2(_07287_),
    .B1(_07348_),
    .C1(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__inv_2 _13058_ (.A(_07362_),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _13059_ (.A(\CPU_Xreg_value_a4[5][0] ),
    .Y(_07363_));
 sky130_fd_sc_hd__nor2_4 _13060_ (.A(_07363_),
    .B(_07285_),
    .Y(_07364_));
 sky130_fd_sc_hd__a211o_4 _13061_ (.A1(_07188_),
    .A2(_07285_),
    .B1(_07274_),
    .C1(_07364_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_4 _13062_ (.A(_06986_),
    .B(_07192_),
    .X(_07365_));
 sky130_fd_sc_hd__nor2_4 _13063_ (.A(_06166_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__buf_2 _13064_ (.A(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__buf_2 _13065_ (.A(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__buf_2 _13066_ (.A(_07158_),
    .X(_07369_));
 sky130_fd_sc_hd__buf_2 _13067_ (.A(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_2 _13068_ (.A(_07367_),
    .X(_07371_));
 sky130_fd_sc_hd__nor2_4 _13069_ (.A(\CPU_Xreg_value_a4[6][31] ),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__a211o_4 _13070_ (.A1(_06984_),
    .A2(_07368_),
    .B1(_07370_),
    .C1(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__inv_2 _13071_ (.A(_07373_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_4 _13072_ (.A(\CPU_Xreg_value_a4[6][30] ),
    .B(_07371_),
    .Y(_07374_));
 sky130_fd_sc_hd__a211o_4 _13073_ (.A1(_06994_),
    .A2(_07368_),
    .B1(_07370_),
    .C1(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__inv_2 _13074_ (.A(_07375_),
    .Y(_00844_));
 sky130_fd_sc_hd__buf_2 _13075_ (.A(_07366_),
    .X(_07376_));
 sky130_fd_sc_hd__buf_2 _13076_ (.A(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__buf_2 _13077_ (.A(_07367_),
    .X(_07378_));
 sky130_fd_sc_hd__nor2_4 _13078_ (.A(\CPU_Xreg_value_a4[6][29] ),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__a211o_4 _13079_ (.A1(_06997_),
    .A2(_07377_),
    .B1(_07370_),
    .C1(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__inv_2 _13080_ (.A(_07380_),
    .Y(_00843_));
 sky130_fd_sc_hd__nor2_4 _13081_ (.A(\CPU_Xreg_value_a4[6][28] ),
    .B(_07378_),
    .Y(_07381_));
 sky130_fd_sc_hd__a211o_4 _13082_ (.A1(_07001_),
    .A2(_07377_),
    .B1(_07370_),
    .C1(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__inv_2 _13083_ (.A(_07382_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_4 _13084_ (.A(\CPU_Xreg_value_a4[6][27] ),
    .B(_07378_),
    .Y(_07383_));
 sky130_fd_sc_hd__a211o_4 _13085_ (.A1(_07005_),
    .A2(_07377_),
    .B1(_07370_),
    .C1(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__inv_2 _13086_ (.A(_07384_),
    .Y(_00841_));
 sky130_fd_sc_hd__nor2_4 _13087_ (.A(\CPU_Xreg_value_a4[6][26] ),
    .B(_07378_),
    .Y(_07385_));
 sky130_fd_sc_hd__a211o_4 _13088_ (.A1(_07010_),
    .A2(_07377_),
    .B1(_07370_),
    .C1(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__inv_2 _13089_ (.A(_07386_),
    .Y(_00840_));
 sky130_fd_sc_hd__buf_2 _13090_ (.A(_07369_),
    .X(_07387_));
 sky130_fd_sc_hd__nor2_4 _13091_ (.A(\CPU_Xreg_value_a4[6][25] ),
    .B(_07378_),
    .Y(_07388_));
 sky130_fd_sc_hd__a211o_4 _13092_ (.A1(_07013_),
    .A2(_07377_),
    .B1(_07387_),
    .C1(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__inv_2 _13093_ (.A(_07389_),
    .Y(_00839_));
 sky130_fd_sc_hd__nor2_4 _13094_ (.A(\CPU_Xreg_value_a4[6][24] ),
    .B(_07378_),
    .Y(_07390_));
 sky130_fd_sc_hd__a211o_4 _13095_ (.A1(_07016_),
    .A2(_07377_),
    .B1(_07387_),
    .C1(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__inv_2 _13096_ (.A(_07391_),
    .Y(_00838_));
 sky130_fd_sc_hd__buf_2 _13097_ (.A(_07376_),
    .X(_07392_));
 sky130_fd_sc_hd__buf_2 _13098_ (.A(_07367_),
    .X(_07393_));
 sky130_fd_sc_hd__nor2_4 _13099_ (.A(\CPU_Xreg_value_a4[6][23] ),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__a211o_4 _13100_ (.A1(_07019_),
    .A2(_07392_),
    .B1(_07387_),
    .C1(_07394_),
    .X(_07395_));
 sky130_fd_sc_hd__inv_2 _13101_ (.A(_07395_),
    .Y(_00837_));
 sky130_fd_sc_hd__nor2_4 _13102_ (.A(\CPU_Xreg_value_a4[6][22] ),
    .B(_07393_),
    .Y(_07396_));
 sky130_fd_sc_hd__a211o_4 _13103_ (.A1(_07023_),
    .A2(_07392_),
    .B1(_07387_),
    .C1(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__inv_2 _13104_ (.A(_07397_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2_4 _13105_ (.A(\CPU_Xreg_value_a4[6][21] ),
    .B(_07393_),
    .Y(_07398_));
 sky130_fd_sc_hd__a211o_4 _13106_ (.A1(_07027_),
    .A2(_07392_),
    .B1(_07387_),
    .C1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__inv_2 _13107_ (.A(_07399_),
    .Y(_00835_));
 sky130_fd_sc_hd__nor2_4 _13108_ (.A(\CPU_Xreg_value_a4[6][20] ),
    .B(_07393_),
    .Y(_07400_));
 sky130_fd_sc_hd__a211o_4 _13109_ (.A1(_07031_),
    .A2(_07392_),
    .B1(_07387_),
    .C1(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(_07401_),
    .Y(_00834_));
 sky130_fd_sc_hd__buf_2 _13111_ (.A(_07369_),
    .X(_07402_));
 sky130_fd_sc_hd__nor2_4 _13112_ (.A(\CPU_Xreg_value_a4[6][19] ),
    .B(_07393_),
    .Y(_07403_));
 sky130_fd_sc_hd__a211o_4 _13113_ (.A1(_07034_),
    .A2(_07392_),
    .B1(_07402_),
    .C1(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__inv_2 _13114_ (.A(_07404_),
    .Y(_00833_));
 sky130_fd_sc_hd__nor2_4 _13115_ (.A(\CPU_Xreg_value_a4[6][18] ),
    .B(_07393_),
    .Y(_07405_));
 sky130_fd_sc_hd__a211o_4 _13116_ (.A1(_07037_),
    .A2(_07392_),
    .B1(_07402_),
    .C1(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__inv_2 _13117_ (.A(_07406_),
    .Y(_00832_));
 sky130_fd_sc_hd__buf_2 _13118_ (.A(_07367_),
    .X(_07407_));
 sky130_fd_sc_hd__buf_2 _13119_ (.A(_07366_),
    .X(_07408_));
 sky130_fd_sc_hd__nor2_4 _13120_ (.A(\CPU_Xreg_value_a4[6][17] ),
    .B(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__a211o_4 _13121_ (.A1(_07040_),
    .A2(_07407_),
    .B1(_07402_),
    .C1(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__inv_2 _13122_ (.A(_07410_),
    .Y(_00831_));
 sky130_fd_sc_hd__nor2_4 _13123_ (.A(\CPU_Xreg_value_a4[6][16] ),
    .B(_07408_),
    .Y(_07411_));
 sky130_fd_sc_hd__a211o_4 _13124_ (.A1(_07045_),
    .A2(_07407_),
    .B1(_07402_),
    .C1(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__inv_2 _13125_ (.A(_07412_),
    .Y(_00830_));
 sky130_fd_sc_hd__nor2_4 _13126_ (.A(\CPU_Xreg_value_a4[6][15] ),
    .B(_07408_),
    .Y(_07413_));
 sky130_fd_sc_hd__a211o_4 _13127_ (.A1(_07049_),
    .A2(_07407_),
    .B1(_07402_),
    .C1(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__inv_2 _13128_ (.A(_07414_),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_4 _13129_ (.A(\CPU_Xreg_value_a4[6][14] ),
    .B(_07408_),
    .Y(_07415_));
 sky130_fd_sc_hd__a211o_4 _13130_ (.A1(_07053_),
    .A2(_07407_),
    .B1(_07402_),
    .C1(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__inv_2 _13131_ (.A(_07416_),
    .Y(_00828_));
 sky130_fd_sc_hd__buf_2 _13132_ (.A(_07369_),
    .X(_07417_));
 sky130_fd_sc_hd__nor2_4 _13133_ (.A(\CPU_Xreg_value_a4[6][13] ),
    .B(_07408_),
    .Y(_07418_));
 sky130_fd_sc_hd__a211o_4 _13134_ (.A1(_07056_),
    .A2(_07407_),
    .B1(_07417_),
    .C1(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__inv_2 _13135_ (.A(_07419_),
    .Y(_00827_));
 sky130_fd_sc_hd__nor2_4 _13136_ (.A(\CPU_Xreg_value_a4[6][12] ),
    .B(_07408_),
    .Y(_07420_));
 sky130_fd_sc_hd__a211o_4 _13137_ (.A1(_07059_),
    .A2(_07407_),
    .B1(_07417_),
    .C1(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__inv_2 _13138_ (.A(_07421_),
    .Y(_00826_));
 sky130_fd_sc_hd__buf_2 _13139_ (.A(_07367_),
    .X(_07422_));
 sky130_fd_sc_hd__buf_2 _13140_ (.A(_07366_),
    .X(_07423_));
 sky130_fd_sc_hd__nor2_4 _13141_ (.A(\CPU_Xreg_value_a4[6][11] ),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__a211o_4 _13142_ (.A1(_07062_),
    .A2(_07422_),
    .B1(_07417_),
    .C1(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__inv_2 _13143_ (.A(_07425_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_4 _13144_ (.A(\CPU_Xreg_value_a4[6][10] ),
    .B(_07423_),
    .Y(_07426_));
 sky130_fd_sc_hd__a211o_4 _13145_ (.A1(_07066_),
    .A2(_07422_),
    .B1(_07417_),
    .C1(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__inv_2 _13146_ (.A(_07427_),
    .Y(_00824_));
 sky130_fd_sc_hd__nor2_4 _13147_ (.A(\CPU_Xreg_value_a4[6][9] ),
    .B(_07423_),
    .Y(_07428_));
 sky130_fd_sc_hd__a211o_4 _13148_ (.A1(_07070_),
    .A2(_07422_),
    .B1(_07417_),
    .C1(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__inv_2 _13149_ (.A(_07429_),
    .Y(_00823_));
 sky130_fd_sc_hd__nor2_4 _13150_ (.A(\CPU_Xreg_value_a4[6][8] ),
    .B(_07423_),
    .Y(_07430_));
 sky130_fd_sc_hd__a211o_4 _13151_ (.A1(_07074_),
    .A2(_07422_),
    .B1(_07417_),
    .C1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__inv_2 _13152_ (.A(_07431_),
    .Y(_00822_));
 sky130_fd_sc_hd__buf_2 _13153_ (.A(_07369_),
    .X(_07432_));
 sky130_fd_sc_hd__nor2_4 _13154_ (.A(\CPU_Xreg_value_a4[6][7] ),
    .B(_07423_),
    .Y(_07433_));
 sky130_fd_sc_hd__a211o_4 _13155_ (.A1(_07077_),
    .A2(_07422_),
    .B1(_07432_),
    .C1(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__inv_2 _13156_ (.A(_07434_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_4 _13157_ (.A(\CPU_Xreg_value_a4[6][6] ),
    .B(_07423_),
    .Y(_07435_));
 sky130_fd_sc_hd__a211o_4 _13158_ (.A1(_07080_),
    .A2(_07422_),
    .B1(_07432_),
    .C1(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__inv_2 _13159_ (.A(_07436_),
    .Y(_00820_));
 sky130_fd_sc_hd__nor2_4 _13160_ (.A(\CPU_Xreg_value_a4[6][5] ),
    .B(_07376_),
    .Y(_07437_));
 sky130_fd_sc_hd__a211o_4 _13161_ (.A1(_07083_),
    .A2(_07371_),
    .B1(_07432_),
    .C1(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__inv_2 _13162_ (.A(_07438_),
    .Y(_00819_));
 sky130_fd_sc_hd__nor2_4 _13163_ (.A(\CPU_Xreg_value_a4[6][4] ),
    .B(_07376_),
    .Y(_07439_));
 sky130_fd_sc_hd__a211o_4 _13164_ (.A1(_07087_),
    .A2(_07371_),
    .B1(_07432_),
    .C1(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__inv_2 _13165_ (.A(_07440_),
    .Y(_00818_));
 sky130_fd_sc_hd__nor2_4 _13166_ (.A(\CPU_Xreg_value_a4[6][3] ),
    .B(_07376_),
    .Y(_07441_));
 sky130_fd_sc_hd__a211o_4 _13167_ (.A1(_07090_),
    .A2(_07371_),
    .B1(_07432_),
    .C1(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__inv_2 _13168_ (.A(_07442_),
    .Y(_00817_));
 sky130_fd_sc_hd__inv_2 _13169_ (.A(\CPU_Xreg_value_a4[6][2] ),
    .Y(_07443_));
 sky130_fd_sc_hd__nor2_4 _13170_ (.A(_07443_),
    .B(_07368_),
    .Y(_07444_));
 sky130_fd_sc_hd__a211o_4 _13171_ (.A1(_07272_),
    .A2(_07368_),
    .B1(_07274_),
    .C1(_07444_),
    .X(_00816_));
 sky130_fd_sc_hd__inv_2 _13172_ (.A(\CPU_Xreg_value_a4[6][1] ),
    .Y(_07445_));
 sky130_fd_sc_hd__nor2_4 _13173_ (.A(_07445_),
    .B(_07368_),
    .Y(_07446_));
 sky130_fd_sc_hd__a211o_4 _13174_ (.A1(_07097_),
    .A2(_07368_),
    .B1(_07274_),
    .C1(_07446_),
    .X(_00815_));
 sky130_fd_sc_hd__nor2_4 _13175_ (.A(\CPU_Xreg_value_a4[6][0] ),
    .B(_07376_),
    .Y(_07447_));
 sky130_fd_sc_hd__a211o_4 _13176_ (.A1(_07101_),
    .A2(_07371_),
    .B1(_07432_),
    .C1(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__inv_2 _13177_ (.A(_07448_),
    .Y(_00814_));
 sky130_fd_sc_hd__buf_2 _13178_ (.A(_06165_),
    .X(_07449_));
 sky130_fd_sc_hd__or2_4 _13179_ (.A(_07104_),
    .B(_07192_),
    .X(_07450_));
 sky130_fd_sc_hd__nor2_4 _13180_ (.A(_07449_),
    .B(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__buf_2 _13181_ (.A(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__buf_2 _13182_ (.A(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__buf_2 _13183_ (.A(_07369_),
    .X(_07454_));
 sky130_fd_sc_hd__buf_2 _13184_ (.A(_07451_),
    .X(_07455_));
 sky130_fd_sc_hd__buf_2 _13185_ (.A(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__nor2_4 _13186_ (.A(\CPU_Xreg_value_a4[7][31] ),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__a211o_4 _13187_ (.A1(_06984_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__inv_2 _13188_ (.A(_07458_),
    .Y(_00813_));
 sky130_fd_sc_hd__buf_2 _13189_ (.A(_07455_),
    .X(_07459_));
 sky130_fd_sc_hd__nor2_4 _13190_ (.A(\CPU_Xreg_value_a4[7][30] ),
    .B(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__a211o_4 _13191_ (.A1(_06994_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07460_),
    .X(_07461_));
 sky130_fd_sc_hd__inv_2 _13192_ (.A(_07461_),
    .Y(_00812_));
 sky130_fd_sc_hd__nor2_4 _13193_ (.A(\CPU_Xreg_value_a4[7][29] ),
    .B(_07459_),
    .Y(_07462_));
 sky130_fd_sc_hd__a211o_4 _13194_ (.A1(_06997_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__inv_2 _13195_ (.A(_07463_),
    .Y(_00811_));
 sky130_fd_sc_hd__nor2_4 _13196_ (.A(\CPU_Xreg_value_a4[7][28] ),
    .B(_07459_),
    .Y(_07464_));
 sky130_fd_sc_hd__a211o_4 _13197_ (.A1(_07001_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__inv_2 _13198_ (.A(_07465_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor2_4 _13199_ (.A(\CPU_Xreg_value_a4[7][27] ),
    .B(_07459_),
    .Y(_07466_));
 sky130_fd_sc_hd__a211o_4 _13200_ (.A1(_07005_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__inv_2 _13201_ (.A(_07467_),
    .Y(_00809_));
 sky130_fd_sc_hd__nor2_4 _13202_ (.A(\CPU_Xreg_value_a4[7][26] ),
    .B(_07459_),
    .Y(_07468_));
 sky130_fd_sc_hd__a211o_4 _13203_ (.A1(_07010_),
    .A2(_07453_),
    .B1(_07454_),
    .C1(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__inv_2 _13204_ (.A(_07469_),
    .Y(_00808_));
 sky130_fd_sc_hd__buf_2 _13205_ (.A(_07455_),
    .X(_07470_));
 sky130_fd_sc_hd__buf_2 _13206_ (.A(_07158_),
    .X(_07471_));
 sky130_fd_sc_hd__buf_2 _13207_ (.A(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__nor2_4 _13208_ (.A(\CPU_Xreg_value_a4[7][25] ),
    .B(_07459_),
    .Y(_07473_));
 sky130_fd_sc_hd__a211o_4 _13209_ (.A1(_07013_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07473_),
    .X(_07474_));
 sky130_fd_sc_hd__inv_2 _13210_ (.A(_07474_),
    .Y(_00807_));
 sky130_fd_sc_hd__buf_2 _13211_ (.A(_07455_),
    .X(_07475_));
 sky130_fd_sc_hd__nor2_4 _13212_ (.A(\CPU_Xreg_value_a4[7][24] ),
    .B(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__a211o_4 _13213_ (.A1(_07016_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__inv_2 _13214_ (.A(_07477_),
    .Y(_00806_));
 sky130_fd_sc_hd__nor2_4 _13215_ (.A(\CPU_Xreg_value_a4[7][23] ),
    .B(_07475_),
    .Y(_07478_));
 sky130_fd_sc_hd__a211o_4 _13216_ (.A1(_07019_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07478_),
    .X(_07479_));
 sky130_fd_sc_hd__inv_2 _13217_ (.A(_07479_),
    .Y(_00805_));
 sky130_fd_sc_hd__nor2_4 _13218_ (.A(\CPU_Xreg_value_a4[7][22] ),
    .B(_07475_),
    .Y(_07480_));
 sky130_fd_sc_hd__a211o_4 _13219_ (.A1(_07023_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__inv_2 _13220_ (.A(_07481_),
    .Y(_00804_));
 sky130_fd_sc_hd__nor2_4 _13221_ (.A(\CPU_Xreg_value_a4[7][21] ),
    .B(_07475_),
    .Y(_07482_));
 sky130_fd_sc_hd__a211o_4 _13222_ (.A1(_07027_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__inv_2 _13223_ (.A(_07483_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_4 _13224_ (.A(\CPU_Xreg_value_a4[7][20] ),
    .B(_07475_),
    .Y(_07484_));
 sky130_fd_sc_hd__a211o_4 _13225_ (.A1(_07031_),
    .A2(_07470_),
    .B1(_07472_),
    .C1(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__inv_2 _13226_ (.A(_07485_),
    .Y(_00802_));
 sky130_fd_sc_hd__buf_2 _13227_ (.A(_07455_),
    .X(_07486_));
 sky130_fd_sc_hd__buf_2 _13228_ (.A(_07471_),
    .X(_07487_));
 sky130_fd_sc_hd__nor2_4 _13229_ (.A(\CPU_Xreg_value_a4[7][19] ),
    .B(_07475_),
    .Y(_07488_));
 sky130_fd_sc_hd__a211o_4 _13230_ (.A1(_07034_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__inv_2 _13231_ (.A(_07489_),
    .Y(_00801_));
 sky130_fd_sc_hd__buf_2 _13232_ (.A(_07451_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_4 _13233_ (.A(\CPU_Xreg_value_a4[7][18] ),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__a211o_4 _13234_ (.A1(_07037_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__inv_2 _13235_ (.A(_07492_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor2_4 _13236_ (.A(\CPU_Xreg_value_a4[7][17] ),
    .B(_07490_),
    .Y(_07493_));
 sky130_fd_sc_hd__a211o_4 _13237_ (.A1(_07040_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__inv_2 _13238_ (.A(_07494_),
    .Y(_00799_));
 sky130_fd_sc_hd__nor2_4 _13239_ (.A(\CPU_Xreg_value_a4[7][16] ),
    .B(_07490_),
    .Y(_07495_));
 sky130_fd_sc_hd__a211o_4 _13240_ (.A1(_07045_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__inv_2 _13241_ (.A(_07496_),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_4 _13242_ (.A(\CPU_Xreg_value_a4[7][15] ),
    .B(_07490_),
    .Y(_07497_));
 sky130_fd_sc_hd__a211o_4 _13243_ (.A1(_07049_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__inv_2 _13244_ (.A(_07498_),
    .Y(_00797_));
 sky130_fd_sc_hd__nor2_4 _13245_ (.A(\CPU_Xreg_value_a4[7][14] ),
    .B(_07490_),
    .Y(_07499_));
 sky130_fd_sc_hd__a211o_4 _13246_ (.A1(_07053_),
    .A2(_07486_),
    .B1(_07487_),
    .C1(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__inv_2 _13247_ (.A(_07500_),
    .Y(_00796_));
 sky130_fd_sc_hd__buf_2 _13248_ (.A(_07455_),
    .X(_07501_));
 sky130_fd_sc_hd__buf_2 _13249_ (.A(_07471_),
    .X(_07502_));
 sky130_fd_sc_hd__nor2_4 _13250_ (.A(\CPU_Xreg_value_a4[7][13] ),
    .B(_07490_),
    .Y(_07503_));
 sky130_fd_sc_hd__a211o_4 _13251_ (.A1(_07056_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__inv_2 _13252_ (.A(_07504_),
    .Y(_00795_));
 sky130_fd_sc_hd__buf_2 _13253_ (.A(_07451_),
    .X(_07505_));
 sky130_fd_sc_hd__nor2_4 _13254_ (.A(\CPU_Xreg_value_a4[7][12] ),
    .B(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__a211o_4 _13255_ (.A1(_07059_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07506_),
    .X(_07507_));
 sky130_fd_sc_hd__inv_2 _13256_ (.A(_07507_),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_4 _13257_ (.A(\CPU_Xreg_value_a4[7][11] ),
    .B(_07505_),
    .Y(_07508_));
 sky130_fd_sc_hd__a211o_4 _13258_ (.A1(_07062_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__inv_2 _13259_ (.A(_07509_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_4 _13260_ (.A(\CPU_Xreg_value_a4[7][10] ),
    .B(_07505_),
    .Y(_07510_));
 sky130_fd_sc_hd__a211o_4 _13261_ (.A1(_07066_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__inv_2 _13262_ (.A(_07511_),
    .Y(_00792_));
 sky130_fd_sc_hd__nor2_4 _13263_ (.A(\CPU_Xreg_value_a4[7][9] ),
    .B(_07505_),
    .Y(_07512_));
 sky130_fd_sc_hd__a211o_4 _13264_ (.A1(_07070_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__inv_2 _13265_ (.A(_07513_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_4 _13266_ (.A(\CPU_Xreg_value_a4[7][8] ),
    .B(_07505_),
    .Y(_07514_));
 sky130_fd_sc_hd__a211o_4 _13267_ (.A1(_07074_),
    .A2(_07501_),
    .B1(_07502_),
    .C1(_07514_),
    .X(_07515_));
 sky130_fd_sc_hd__inv_2 _13268_ (.A(_07515_),
    .Y(_00790_));
 sky130_fd_sc_hd__buf_2 _13269_ (.A(_07471_),
    .X(_07516_));
 sky130_fd_sc_hd__nor2_4 _13270_ (.A(\CPU_Xreg_value_a4[7][7] ),
    .B(_07505_),
    .Y(_07517_));
 sky130_fd_sc_hd__a211o_4 _13271_ (.A1(_07077_),
    .A2(_07456_),
    .B1(_07516_),
    .C1(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__inv_2 _13272_ (.A(_07518_),
    .Y(_00789_));
 sky130_fd_sc_hd__nor2_4 _13273_ (.A(\CPU_Xreg_value_a4[7][6] ),
    .B(_07452_),
    .Y(_07519_));
 sky130_fd_sc_hd__a211o_4 _13274_ (.A1(_07080_),
    .A2(_07456_),
    .B1(_07516_),
    .C1(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__inv_2 _13275_ (.A(_07520_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor2_4 _13276_ (.A(\CPU_Xreg_value_a4[7][5] ),
    .B(_07452_),
    .Y(_07521_));
 sky130_fd_sc_hd__a211o_4 _13277_ (.A1(_07083_),
    .A2(_07456_),
    .B1(_07516_),
    .C1(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__inv_2 _13278_ (.A(_07522_),
    .Y(_00787_));
 sky130_fd_sc_hd__nor2_4 _13279_ (.A(\CPU_Xreg_value_a4[7][4] ),
    .B(_07452_),
    .Y(_07523_));
 sky130_fd_sc_hd__a211o_4 _13280_ (.A1(_07087_),
    .A2(_07456_),
    .B1(_07516_),
    .C1(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__inv_2 _13281_ (.A(_07524_),
    .Y(_00786_));
 sky130_fd_sc_hd__nor2_4 _13282_ (.A(\CPU_Xreg_value_a4[7][3] ),
    .B(_07452_),
    .Y(_07525_));
 sky130_fd_sc_hd__a211o_4 _13283_ (.A1(_07090_),
    .A2(_07456_),
    .B1(_07516_),
    .C1(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__inv_2 _13284_ (.A(_07526_),
    .Y(_00785_));
 sky130_fd_sc_hd__buf_2 _13285_ (.A(_07452_),
    .X(_07527_));
 sky130_fd_sc_hd__inv_2 _13286_ (.A(\CPU_Xreg_value_a4[7][2] ),
    .Y(_07528_));
 sky130_fd_sc_hd__nor2_4 _13287_ (.A(_07528_),
    .B(_07527_),
    .Y(_07529_));
 sky130_fd_sc_hd__a211o_4 _13288_ (.A1(_07272_),
    .A2(_07527_),
    .B1(_07274_),
    .C1(_07529_),
    .X(_00784_));
 sky130_fd_sc_hd__buf_2 _13289_ (.A(_07273_),
    .X(_07530_));
 sky130_fd_sc_hd__inv_2 _13290_ (.A(\CPU_Xreg_value_a4[7][1] ),
    .Y(_07531_));
 sky130_fd_sc_hd__nor2_4 _13291_ (.A(_07531_),
    .B(_07527_),
    .Y(_07532_));
 sky130_fd_sc_hd__a211o_4 _13292_ (.A1(_07097_),
    .A2(_07527_),
    .B1(_07530_),
    .C1(_07532_),
    .X(_00783_));
 sky130_fd_sc_hd__inv_2 _13293_ (.A(\CPU_Xreg_value_a4[7][0] ),
    .Y(_07533_));
 sky130_fd_sc_hd__nor2_4 _13294_ (.A(_07533_),
    .B(_07527_),
    .Y(_07534_));
 sky130_fd_sc_hd__a211o_4 _13295_ (.A1(_07188_),
    .A2(_07527_),
    .B1(_07530_),
    .C1(_07534_),
    .X(_00782_));
 sky130_fd_sc_hd__buf_2 _13296_ (.A(_06503_),
    .X(_07535_));
 sky130_fd_sc_hd__inv_2 _13297_ (.A(_06147_),
    .Y(_07536_));
 sky130_fd_sc_hd__or2_4 _13298_ (.A(_06145_),
    .B(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__or2_4 _13299_ (.A(_06156_),
    .B(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__nor2_4 _13300_ (.A(_07449_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__buf_2 _13301_ (.A(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__buf_2 _13302_ (.A(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__buf_2 _13303_ (.A(_07540_),
    .X(_07542_));
 sky130_fd_sc_hd__nor2_4 _13304_ (.A(\CPU_Xreg_value_a4[8][31] ),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__a211o_4 _13305_ (.A1(_07535_),
    .A2(_07541_),
    .B1(_07516_),
    .C1(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__inv_2 _13306_ (.A(_07544_),
    .Y(_00781_));
 sky130_fd_sc_hd__buf_2 _13307_ (.A(_06515_),
    .X(_07545_));
 sky130_fd_sc_hd__buf_2 _13308_ (.A(_07471_),
    .X(_07546_));
 sky130_fd_sc_hd__nor2_4 _13309_ (.A(\CPU_Xreg_value_a4[8][30] ),
    .B(_07542_),
    .Y(_07547_));
 sky130_fd_sc_hd__a211o_4 _13310_ (.A1(_07545_),
    .A2(_07541_),
    .B1(_07546_),
    .C1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__inv_2 _13311_ (.A(_07548_),
    .Y(_00780_));
 sky130_fd_sc_hd__buf_2 _13312_ (.A(_06531_),
    .X(_07549_));
 sky130_fd_sc_hd__nor2_4 _13313_ (.A(\CPU_Xreg_value_a4[8][29] ),
    .B(_07542_),
    .Y(_07550_));
 sky130_fd_sc_hd__a211o_4 _13314_ (.A1(_07549_),
    .A2(_07541_),
    .B1(_07546_),
    .C1(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__inv_2 _13315_ (.A(_07551_),
    .Y(_00779_));
 sky130_fd_sc_hd__buf_2 _13316_ (.A(_06539_),
    .X(_07552_));
 sky130_fd_sc_hd__buf_2 _13317_ (.A(_07540_),
    .X(_07553_));
 sky130_fd_sc_hd__nor2_4 _13318_ (.A(\CPU_Xreg_value_a4[8][28] ),
    .B(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__a211o_4 _13319_ (.A1(_07552_),
    .A2(_07541_),
    .B1(_07546_),
    .C1(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__inv_2 _13320_ (.A(_07555_),
    .Y(_00778_));
 sky130_fd_sc_hd__buf_2 _13321_ (.A(_06564_),
    .X(_07556_));
 sky130_fd_sc_hd__buf_2 _13322_ (.A(_07539_),
    .X(_07557_));
 sky130_fd_sc_hd__buf_2 _13323_ (.A(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__nor2_4 _13324_ (.A(\CPU_Xreg_value_a4[8][27] ),
    .B(_07553_),
    .Y(_07559_));
 sky130_fd_sc_hd__a211o_4 _13325_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_07546_),
    .C1(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__inv_2 _13326_ (.A(_07560_),
    .Y(_00777_));
 sky130_fd_sc_hd__buf_2 _13327_ (.A(_06574_),
    .X(_07561_));
 sky130_fd_sc_hd__nor2_4 _13328_ (.A(\CPU_Xreg_value_a4[8][26] ),
    .B(_07553_),
    .Y(_07562_));
 sky130_fd_sc_hd__a211o_4 _13329_ (.A1(_07561_),
    .A2(_07558_),
    .B1(_07546_),
    .C1(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__inv_2 _13330_ (.A(_07563_),
    .Y(_00776_));
 sky130_fd_sc_hd__buf_2 _13331_ (.A(_06589_),
    .X(_07564_));
 sky130_fd_sc_hd__nor2_4 _13332_ (.A(\CPU_Xreg_value_a4[8][25] ),
    .B(_07553_),
    .Y(_07565_));
 sky130_fd_sc_hd__a211o_4 _13333_ (.A1(_07564_),
    .A2(_07558_),
    .B1(_07546_),
    .C1(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__inv_2 _13334_ (.A(_07566_),
    .Y(_00775_));
 sky130_fd_sc_hd__buf_2 _13335_ (.A(_06599_),
    .X(_07567_));
 sky130_fd_sc_hd__buf_2 _13336_ (.A(_07471_),
    .X(_07568_));
 sky130_fd_sc_hd__nor2_4 _13337_ (.A(\CPU_Xreg_value_a4[8][24] ),
    .B(_07553_),
    .Y(_07569_));
 sky130_fd_sc_hd__a211o_4 _13338_ (.A1(_07567_),
    .A2(_07558_),
    .B1(_07568_),
    .C1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__inv_2 _13339_ (.A(_07570_),
    .Y(_00774_));
 sky130_fd_sc_hd__buf_2 _13340_ (.A(_06619_),
    .X(_07571_));
 sky130_fd_sc_hd__nor2_4 _13341_ (.A(\CPU_Xreg_value_a4[8][23] ),
    .B(_07553_),
    .Y(_07572_));
 sky130_fd_sc_hd__a211o_4 _13342_ (.A1(_07571_),
    .A2(_07558_),
    .B1(_07568_),
    .C1(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__inv_2 _13343_ (.A(_07573_),
    .Y(_00773_));
 sky130_fd_sc_hd__buf_2 _13344_ (.A(_06627_),
    .X(_07574_));
 sky130_fd_sc_hd__buf_2 _13345_ (.A(_07540_),
    .X(_07575_));
 sky130_fd_sc_hd__nor2_4 _13346_ (.A(\CPU_Xreg_value_a4[8][22] ),
    .B(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__a211o_4 _13347_ (.A1(_07574_),
    .A2(_07558_),
    .B1(_07568_),
    .C1(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__inv_2 _13348_ (.A(_07577_),
    .Y(_00772_));
 sky130_fd_sc_hd__buf_2 _13349_ (.A(_06642_),
    .X(_07578_));
 sky130_fd_sc_hd__buf_2 _13350_ (.A(_07557_),
    .X(_07579_));
 sky130_fd_sc_hd__nor2_4 _13351_ (.A(\CPU_Xreg_value_a4[8][21] ),
    .B(_07575_),
    .Y(_07580_));
 sky130_fd_sc_hd__a211o_4 _13352_ (.A1(_07578_),
    .A2(_07579_),
    .B1(_07568_),
    .C1(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__inv_2 _13353_ (.A(_07581_),
    .Y(_00771_));
 sky130_fd_sc_hd__buf_2 _13354_ (.A(_06651_),
    .X(_07582_));
 sky130_fd_sc_hd__nor2_4 _13355_ (.A(\CPU_Xreg_value_a4[8][20] ),
    .B(_07575_),
    .Y(_07583_));
 sky130_fd_sc_hd__a211o_4 _13356_ (.A1(_07582_),
    .A2(_07579_),
    .B1(_07568_),
    .C1(_07583_),
    .X(_07584_));
 sky130_fd_sc_hd__inv_2 _13357_ (.A(_07584_),
    .Y(_00770_));
 sky130_fd_sc_hd__buf_2 _13358_ (.A(_06673_),
    .X(_07585_));
 sky130_fd_sc_hd__nor2_4 _13359_ (.A(\CPU_Xreg_value_a4[8][19] ),
    .B(_07575_),
    .Y(_07586_));
 sky130_fd_sc_hd__a211o_4 _13360_ (.A1(_07585_),
    .A2(_07579_),
    .B1(_07568_),
    .C1(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__inv_2 _13361_ (.A(_07587_),
    .Y(_00769_));
 sky130_fd_sc_hd__buf_2 _13362_ (.A(_06682_),
    .X(_07588_));
 sky130_fd_sc_hd__buf_2 _13363_ (.A(_07158_),
    .X(_07589_));
 sky130_fd_sc_hd__buf_2 _13364_ (.A(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__nor2_4 _13365_ (.A(\CPU_Xreg_value_a4[8][18] ),
    .B(_07575_),
    .Y(_07591_));
 sky130_fd_sc_hd__a211o_4 _13366_ (.A1(_07588_),
    .A2(_07579_),
    .B1(_07590_),
    .C1(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__inv_2 _13367_ (.A(_07592_),
    .Y(_00768_));
 sky130_fd_sc_hd__buf_2 _13368_ (.A(_06692_),
    .X(_07593_));
 sky130_fd_sc_hd__nor2_4 _13369_ (.A(\CPU_Xreg_value_a4[8][17] ),
    .B(_07575_),
    .Y(_07594_));
 sky130_fd_sc_hd__a211o_4 _13370_ (.A1(_07593_),
    .A2(_07579_),
    .B1(_07590_),
    .C1(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__inv_2 _13371_ (.A(_07595_),
    .Y(_00767_));
 sky130_fd_sc_hd__buf_2 _13372_ (.A(_06701_),
    .X(_07596_));
 sky130_fd_sc_hd__buf_2 _13373_ (.A(_07539_),
    .X(_07597_));
 sky130_fd_sc_hd__nor2_4 _13374_ (.A(\CPU_Xreg_value_a4[8][16] ),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__a211o_4 _13375_ (.A1(_07596_),
    .A2(_07579_),
    .B1(_07590_),
    .C1(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__inv_2 _13376_ (.A(_07599_),
    .Y(_00766_));
 sky130_fd_sc_hd__buf_2 _13377_ (.A(_06724_),
    .X(_07600_));
 sky130_fd_sc_hd__buf_2 _13378_ (.A(_07540_),
    .X(_07601_));
 sky130_fd_sc_hd__nor2_4 _13379_ (.A(\CPU_Xreg_value_a4[8][15] ),
    .B(_07597_),
    .Y(_07602_));
 sky130_fd_sc_hd__a211o_4 _13380_ (.A1(_07600_),
    .A2(_07601_),
    .B1(_07590_),
    .C1(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__inv_2 _13381_ (.A(_07603_),
    .Y(_00765_));
 sky130_fd_sc_hd__buf_2 _13382_ (.A(_06733_),
    .X(_07604_));
 sky130_fd_sc_hd__nor2_4 _13383_ (.A(\CPU_Xreg_value_a4[8][14] ),
    .B(_07597_),
    .Y(_07605_));
 sky130_fd_sc_hd__a211o_4 _13384_ (.A1(_07604_),
    .A2(_07601_),
    .B1(_07590_),
    .C1(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__inv_2 _13385_ (.A(_07606_),
    .Y(_00764_));
 sky130_fd_sc_hd__buf_2 _13386_ (.A(_06743_),
    .X(_07607_));
 sky130_fd_sc_hd__nor2_4 _13387_ (.A(\CPU_Xreg_value_a4[8][13] ),
    .B(_07597_),
    .Y(_07608_));
 sky130_fd_sc_hd__a211o_4 _13388_ (.A1(_07607_),
    .A2(_07601_),
    .B1(_07590_),
    .C1(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__inv_2 _13389_ (.A(_07609_),
    .Y(_00763_));
 sky130_fd_sc_hd__buf_2 _13390_ (.A(_06752_),
    .X(_07610_));
 sky130_fd_sc_hd__buf_2 _13391_ (.A(_07589_),
    .X(_07611_));
 sky130_fd_sc_hd__nor2_4 _13392_ (.A(\CPU_Xreg_value_a4[8][12] ),
    .B(_07597_),
    .Y(_07612_));
 sky130_fd_sc_hd__a211o_4 _13393_ (.A1(_07610_),
    .A2(_07601_),
    .B1(_07611_),
    .C1(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__inv_2 _13394_ (.A(_07613_),
    .Y(_00762_));
 sky130_fd_sc_hd__buf_2 _13395_ (.A(_06770_),
    .X(_07614_));
 sky130_fd_sc_hd__nor2_4 _13396_ (.A(\CPU_Xreg_value_a4[8][11] ),
    .B(_07597_),
    .Y(_07615_));
 sky130_fd_sc_hd__a211o_4 _13397_ (.A1(_07614_),
    .A2(_07601_),
    .B1(_07611_),
    .C1(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__inv_2 _13398_ (.A(_07616_),
    .Y(_00761_));
 sky130_fd_sc_hd__buf_2 _13399_ (.A(_06778_),
    .X(_07617_));
 sky130_fd_sc_hd__buf_2 _13400_ (.A(_07539_),
    .X(_07618_));
 sky130_fd_sc_hd__nor2_4 _13401_ (.A(\CPU_Xreg_value_a4[8][10] ),
    .B(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__a211o_4 _13402_ (.A1(_07617_),
    .A2(_07601_),
    .B1(_07611_),
    .C1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__inv_2 _13403_ (.A(_07620_),
    .Y(_00760_));
 sky130_fd_sc_hd__buf_2 _13404_ (.A(_06791_),
    .X(_07621_));
 sky130_fd_sc_hd__buf_2 _13405_ (.A(_07540_),
    .X(_07622_));
 sky130_fd_sc_hd__nor2_4 _13406_ (.A(\CPU_Xreg_value_a4[8][9] ),
    .B(_07618_),
    .Y(_07623_));
 sky130_fd_sc_hd__a211o_4 _13407_ (.A1(_07621_),
    .A2(_07622_),
    .B1(_07611_),
    .C1(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__inv_2 _13408_ (.A(_07624_),
    .Y(_00759_));
 sky130_fd_sc_hd__buf_2 _13409_ (.A(_06799_),
    .X(_07625_));
 sky130_fd_sc_hd__nor2_4 _13410_ (.A(\CPU_Xreg_value_a4[8][8] ),
    .B(_07618_),
    .Y(_07626_));
 sky130_fd_sc_hd__a211o_4 _13411_ (.A1(_07625_),
    .A2(_07622_),
    .B1(_07611_),
    .C1(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__inv_2 _13412_ (.A(_07627_),
    .Y(_00758_));
 sky130_fd_sc_hd__buf_2 _13413_ (.A(_06820_),
    .X(_07628_));
 sky130_fd_sc_hd__nor2_4 _13414_ (.A(\CPU_Xreg_value_a4[8][7] ),
    .B(_07618_),
    .Y(_07629_));
 sky130_fd_sc_hd__a211o_4 _13415_ (.A1(_07628_),
    .A2(_07622_),
    .B1(_07611_),
    .C1(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__inv_2 _13416_ (.A(_07630_),
    .Y(_00757_));
 sky130_fd_sc_hd__buf_2 _13417_ (.A(_06828_),
    .X(_07631_));
 sky130_fd_sc_hd__buf_2 _13418_ (.A(_07589_),
    .X(_07632_));
 sky130_fd_sc_hd__nor2_4 _13419_ (.A(\CPU_Xreg_value_a4[8][6] ),
    .B(_07618_),
    .Y(_07633_));
 sky130_fd_sc_hd__a211o_4 _13420_ (.A1(_07631_),
    .A2(_07622_),
    .B1(_07632_),
    .C1(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_07634_),
    .Y(_00756_));
 sky130_fd_sc_hd__buf_2 _13422_ (.A(_06837_),
    .X(_07635_));
 sky130_fd_sc_hd__nor2_4 _13423_ (.A(\CPU_Xreg_value_a4[8][5] ),
    .B(_07618_),
    .Y(_07636_));
 sky130_fd_sc_hd__a211o_4 _13424_ (.A1(_07635_),
    .A2(_07622_),
    .B1(_07632_),
    .C1(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__inv_2 _13425_ (.A(_07637_),
    .Y(_00755_));
 sky130_fd_sc_hd__buf_2 _13426_ (.A(_06843_),
    .X(_07638_));
 sky130_fd_sc_hd__nor2_4 _13427_ (.A(\CPU_Xreg_value_a4[8][4] ),
    .B(_07557_),
    .Y(_07639_));
 sky130_fd_sc_hd__a211o_4 _13428_ (.A1(_07638_),
    .A2(_07622_),
    .B1(_07632_),
    .C1(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__inv_2 _13429_ (.A(_07640_),
    .Y(_00754_));
 sky130_fd_sc_hd__buf_2 _13430_ (.A(_06851_),
    .X(_07641_));
 sky130_fd_sc_hd__buf_2 _13431_ (.A(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__inv_2 _13432_ (.A(\CPU_Xreg_value_a4[8][3] ),
    .Y(_07643_));
 sky130_fd_sc_hd__nor2_4 _13433_ (.A(_07643_),
    .B(_07541_),
    .Y(_07644_));
 sky130_fd_sc_hd__a211o_4 _13434_ (.A1(_07642_),
    .A2(_07541_),
    .B1(_07530_),
    .C1(_07644_),
    .X(_00753_));
 sky130_fd_sc_hd__nor2_4 _13435_ (.A(\CPU_Xreg_value_a4[8][2] ),
    .B(_07557_),
    .Y(_07645_));
 sky130_fd_sc_hd__a211o_4 _13436_ (.A1(_07093_),
    .A2(_07542_),
    .B1(_07632_),
    .C1(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__inv_2 _13437_ (.A(_07646_),
    .Y(_00752_));
 sky130_fd_sc_hd__nor2_4 _13438_ (.A(\CPU_Xreg_value_a4[8][1] ),
    .B(_07557_),
    .Y(_07647_));
 sky130_fd_sc_hd__a211o_4 _13439_ (.A1(_07277_),
    .A2(_07542_),
    .B1(_07632_),
    .C1(_07647_),
    .X(_07648_));
 sky130_fd_sc_hd__inv_2 _13440_ (.A(_07648_),
    .Y(_00751_));
 sky130_fd_sc_hd__nor2_4 _13441_ (.A(\CPU_Xreg_value_a4[8][0] ),
    .B(_07557_),
    .Y(_07649_));
 sky130_fd_sc_hd__a211o_4 _13442_ (.A1(_07101_),
    .A2(_07542_),
    .B1(_07632_),
    .C1(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__inv_2 _13443_ (.A(_07650_),
    .Y(_00750_));
 sky130_fd_sc_hd__or2_4 _13444_ (.A(_06152_),
    .B(_07537_),
    .X(_07651_));
 sky130_fd_sc_hd__nor2_4 _13445_ (.A(_07449_),
    .B(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__buf_2 _13446_ (.A(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__buf_2 _13447_ (.A(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__buf_2 _13448_ (.A(_07589_),
    .X(_07655_));
 sky130_fd_sc_hd__buf_2 _13449_ (.A(_07653_),
    .X(_07656_));
 sky130_fd_sc_hd__nor2_4 _13450_ (.A(\CPU_Xreg_value_a4[9][31] ),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__a211o_4 _13451_ (.A1(_07535_),
    .A2(_07654_),
    .B1(_07655_),
    .C1(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__inv_2 _13452_ (.A(_07658_),
    .Y(_00749_));
 sky130_fd_sc_hd__nor2_4 _13453_ (.A(\CPU_Xreg_value_a4[9][30] ),
    .B(_07656_),
    .Y(_07659_));
 sky130_fd_sc_hd__a211o_4 _13454_ (.A1(_07545_),
    .A2(_07654_),
    .B1(_07655_),
    .C1(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__inv_2 _13455_ (.A(_07660_),
    .Y(_00748_));
 sky130_fd_sc_hd__buf_2 _13456_ (.A(_07652_),
    .X(_07661_));
 sky130_fd_sc_hd__buf_2 _13457_ (.A(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__buf_2 _13458_ (.A(_07653_),
    .X(_07663_));
 sky130_fd_sc_hd__nor2_4 _13459_ (.A(\CPU_Xreg_value_a4[9][29] ),
    .B(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__a211o_4 _13460_ (.A1(_07549_),
    .A2(_07662_),
    .B1(_07655_),
    .C1(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__inv_2 _13461_ (.A(_07665_),
    .Y(_00747_));
 sky130_fd_sc_hd__nor2_4 _13462_ (.A(\CPU_Xreg_value_a4[9][28] ),
    .B(_07663_),
    .Y(_07666_));
 sky130_fd_sc_hd__a211o_4 _13463_ (.A1(_07552_),
    .A2(_07662_),
    .B1(_07655_),
    .C1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__inv_2 _13464_ (.A(_07667_),
    .Y(_00746_));
 sky130_fd_sc_hd__nor2_4 _13465_ (.A(\CPU_Xreg_value_a4[9][27] ),
    .B(_07663_),
    .Y(_07668_));
 sky130_fd_sc_hd__a211o_4 _13466_ (.A1(_07556_),
    .A2(_07662_),
    .B1(_07655_),
    .C1(_07668_),
    .X(_07669_));
 sky130_fd_sc_hd__inv_2 _13467_ (.A(_07669_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor2_4 _13468_ (.A(\CPU_Xreg_value_a4[9][26] ),
    .B(_07663_),
    .Y(_07670_));
 sky130_fd_sc_hd__a211o_4 _13469_ (.A1(_07561_),
    .A2(_07662_),
    .B1(_07655_),
    .C1(_07670_),
    .X(_07671_));
 sky130_fd_sc_hd__inv_2 _13470_ (.A(_07671_),
    .Y(_00744_));
 sky130_fd_sc_hd__buf_2 _13471_ (.A(_07589_),
    .X(_07672_));
 sky130_fd_sc_hd__nor2_4 _13472_ (.A(\CPU_Xreg_value_a4[9][25] ),
    .B(_07663_),
    .Y(_07673_));
 sky130_fd_sc_hd__a211o_4 _13473_ (.A1(_07564_),
    .A2(_07662_),
    .B1(_07672_),
    .C1(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__inv_2 _13474_ (.A(_07674_),
    .Y(_00743_));
 sky130_fd_sc_hd__nor2_4 _13475_ (.A(\CPU_Xreg_value_a4[9][24] ),
    .B(_07663_),
    .Y(_07675_));
 sky130_fd_sc_hd__a211o_4 _13476_ (.A1(_07567_),
    .A2(_07662_),
    .B1(_07672_),
    .C1(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__inv_2 _13477_ (.A(_07676_),
    .Y(_00742_));
 sky130_fd_sc_hd__buf_2 _13478_ (.A(_07661_),
    .X(_07677_));
 sky130_fd_sc_hd__buf_2 _13479_ (.A(_07653_),
    .X(_07678_));
 sky130_fd_sc_hd__nor2_4 _13480_ (.A(\CPU_Xreg_value_a4[9][23] ),
    .B(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__a211o_4 _13481_ (.A1(_07571_),
    .A2(_07677_),
    .B1(_07672_),
    .C1(_07679_),
    .X(_07680_));
 sky130_fd_sc_hd__inv_2 _13482_ (.A(_07680_),
    .Y(_00741_));
 sky130_fd_sc_hd__nor2_4 _13483_ (.A(\CPU_Xreg_value_a4[9][22] ),
    .B(_07678_),
    .Y(_07681_));
 sky130_fd_sc_hd__a211o_4 _13484_ (.A1(_07574_),
    .A2(_07677_),
    .B1(_07672_),
    .C1(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__inv_2 _13485_ (.A(_07682_),
    .Y(_00740_));
 sky130_fd_sc_hd__nor2_4 _13486_ (.A(\CPU_Xreg_value_a4[9][21] ),
    .B(_07678_),
    .Y(_07683_));
 sky130_fd_sc_hd__a211o_4 _13487_ (.A1(_07578_),
    .A2(_07677_),
    .B1(_07672_),
    .C1(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__inv_2 _13488_ (.A(_07684_),
    .Y(_00739_));
 sky130_fd_sc_hd__nor2_4 _13489_ (.A(\CPU_Xreg_value_a4[9][20] ),
    .B(_07678_),
    .Y(_07685_));
 sky130_fd_sc_hd__a211o_4 _13490_ (.A1(_07582_),
    .A2(_07677_),
    .B1(_07672_),
    .C1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__inv_2 _13491_ (.A(_07686_),
    .Y(_00738_));
 sky130_fd_sc_hd__buf_2 _13492_ (.A(_07589_),
    .X(_07687_));
 sky130_fd_sc_hd__nor2_4 _13493_ (.A(\CPU_Xreg_value_a4[9][19] ),
    .B(_07678_),
    .Y(_07688_));
 sky130_fd_sc_hd__a211o_4 _13494_ (.A1(_07585_),
    .A2(_07677_),
    .B1(_07687_),
    .C1(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__inv_2 _13495_ (.A(_07689_),
    .Y(_00737_));
 sky130_fd_sc_hd__nor2_4 _13496_ (.A(\CPU_Xreg_value_a4[9][18] ),
    .B(_07678_),
    .Y(_07690_));
 sky130_fd_sc_hd__a211o_4 _13497_ (.A1(_07588_),
    .A2(_07677_),
    .B1(_07687_),
    .C1(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__inv_2 _13498_ (.A(_07691_),
    .Y(_00736_));
 sky130_fd_sc_hd__buf_2 _13499_ (.A(_07653_),
    .X(_07692_));
 sky130_fd_sc_hd__buf_2 _13500_ (.A(_07652_),
    .X(_07693_));
 sky130_fd_sc_hd__nor2_4 _13501_ (.A(\CPU_Xreg_value_a4[9][17] ),
    .B(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__a211o_4 _13502_ (.A1(_07593_),
    .A2(_07692_),
    .B1(_07687_),
    .C1(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__inv_2 _13503_ (.A(_07695_),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2_4 _13504_ (.A(\CPU_Xreg_value_a4[9][16] ),
    .B(_07693_),
    .Y(_07696_));
 sky130_fd_sc_hd__a211o_4 _13505_ (.A1(_07596_),
    .A2(_07692_),
    .B1(_07687_),
    .C1(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__inv_2 _13506_ (.A(_07697_),
    .Y(_00734_));
 sky130_fd_sc_hd__nor2_4 _13507_ (.A(\CPU_Xreg_value_a4[9][15] ),
    .B(_07693_),
    .Y(_07698_));
 sky130_fd_sc_hd__a211o_4 _13508_ (.A1(_07600_),
    .A2(_07692_),
    .B1(_07687_),
    .C1(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__inv_2 _13509_ (.A(_07699_),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2_4 _13510_ (.A(\CPU_Xreg_value_a4[9][14] ),
    .B(_07693_),
    .Y(_07700_));
 sky130_fd_sc_hd__a211o_4 _13511_ (.A1(_07604_),
    .A2(_07692_),
    .B1(_07687_),
    .C1(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__inv_2 _13512_ (.A(_07701_),
    .Y(_00732_));
 sky130_fd_sc_hd__buf_2 _13513_ (.A(_07158_),
    .X(_07702_));
 sky130_fd_sc_hd__buf_2 _13514_ (.A(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__nor2_4 _13515_ (.A(\CPU_Xreg_value_a4[9][13] ),
    .B(_07693_),
    .Y(_07704_));
 sky130_fd_sc_hd__a211o_4 _13516_ (.A1(_07607_),
    .A2(_07692_),
    .B1(_07703_),
    .C1(_07704_),
    .X(_07705_));
 sky130_fd_sc_hd__inv_2 _13517_ (.A(_07705_),
    .Y(_00731_));
 sky130_fd_sc_hd__nor2_4 _13518_ (.A(\CPU_Xreg_value_a4[9][12] ),
    .B(_07693_),
    .Y(_07706_));
 sky130_fd_sc_hd__a211o_4 _13519_ (.A1(_07610_),
    .A2(_07692_),
    .B1(_07703_),
    .C1(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__inv_2 _13520_ (.A(_07707_),
    .Y(_00730_));
 sky130_fd_sc_hd__buf_2 _13521_ (.A(_07653_),
    .X(_07708_));
 sky130_fd_sc_hd__buf_2 _13522_ (.A(_07652_),
    .X(_07709_));
 sky130_fd_sc_hd__nor2_4 _13523_ (.A(\CPU_Xreg_value_a4[9][11] ),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__a211o_4 _13524_ (.A1(_07614_),
    .A2(_07708_),
    .B1(_07703_),
    .C1(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__inv_2 _13525_ (.A(_07711_),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2_4 _13526_ (.A(\CPU_Xreg_value_a4[9][10] ),
    .B(_07709_),
    .Y(_07712_));
 sky130_fd_sc_hd__a211o_4 _13527_ (.A1(_07617_),
    .A2(_07708_),
    .B1(_07703_),
    .C1(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__inv_2 _13528_ (.A(_07713_),
    .Y(_00728_));
 sky130_fd_sc_hd__nor2_4 _13529_ (.A(\CPU_Xreg_value_a4[9][9] ),
    .B(_07709_),
    .Y(_07714_));
 sky130_fd_sc_hd__a211o_4 _13530_ (.A1(_07621_),
    .A2(_07708_),
    .B1(_07703_),
    .C1(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__inv_2 _13531_ (.A(_07715_),
    .Y(_00727_));
 sky130_fd_sc_hd__nor2_4 _13532_ (.A(\CPU_Xreg_value_a4[9][8] ),
    .B(_07709_),
    .Y(_07716_));
 sky130_fd_sc_hd__a211o_4 _13533_ (.A1(_07625_),
    .A2(_07708_),
    .B1(_07703_),
    .C1(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__inv_2 _13534_ (.A(_07717_),
    .Y(_00726_));
 sky130_fd_sc_hd__buf_2 _13535_ (.A(_07702_),
    .X(_07718_));
 sky130_fd_sc_hd__nor2_4 _13536_ (.A(\CPU_Xreg_value_a4[9][7] ),
    .B(_07709_),
    .Y(_07719_));
 sky130_fd_sc_hd__a211o_4 _13537_ (.A1(_07628_),
    .A2(_07708_),
    .B1(_07718_),
    .C1(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__inv_2 _13538_ (.A(_07720_),
    .Y(_00725_));
 sky130_fd_sc_hd__nor2_4 _13539_ (.A(\CPU_Xreg_value_a4[9][6] ),
    .B(_07709_),
    .Y(_07721_));
 sky130_fd_sc_hd__a211o_4 _13540_ (.A1(_07631_),
    .A2(_07708_),
    .B1(_07718_),
    .C1(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__inv_2 _13541_ (.A(_07722_),
    .Y(_00724_));
 sky130_fd_sc_hd__nor2_4 _13542_ (.A(\CPU_Xreg_value_a4[9][5] ),
    .B(_07661_),
    .Y(_07723_));
 sky130_fd_sc_hd__a211o_4 _13543_ (.A1(_07635_),
    .A2(_07656_),
    .B1(_07718_),
    .C1(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__inv_2 _13544_ (.A(_07724_),
    .Y(_00723_));
 sky130_fd_sc_hd__nor2_4 _13545_ (.A(\CPU_Xreg_value_a4[9][4] ),
    .B(_07661_),
    .Y(_07725_));
 sky130_fd_sc_hd__a211o_4 _13546_ (.A1(_07638_),
    .A2(_07656_),
    .B1(_07718_),
    .C1(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__inv_2 _13547_ (.A(_07726_),
    .Y(_00722_));
 sky130_fd_sc_hd__inv_2 _13548_ (.A(\CPU_Xreg_value_a4[9][3] ),
    .Y(_07727_));
 sky130_fd_sc_hd__nor2_4 _13549_ (.A(_07727_),
    .B(_07654_),
    .Y(_07728_));
 sky130_fd_sc_hd__a211o_4 _13550_ (.A1(_07642_),
    .A2(_07654_),
    .B1(_07530_),
    .C1(_07728_),
    .X(_00721_));
 sky130_fd_sc_hd__nor2_4 _13551_ (.A(\CPU_Xreg_value_a4[9][2] ),
    .B(_07661_),
    .Y(_07729_));
 sky130_fd_sc_hd__a211o_4 _13552_ (.A1(_07093_),
    .A2(_07656_),
    .B1(_07718_),
    .C1(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__inv_2 _13553_ (.A(_07730_),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_4 _13554_ (.A(\CPU_Xreg_value_a4[9][1] ),
    .B(_07661_),
    .Y(_07731_));
 sky130_fd_sc_hd__a211o_4 _13555_ (.A1(_07277_),
    .A2(_07656_),
    .B1(_07718_),
    .C1(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__inv_2 _13556_ (.A(_07732_),
    .Y(_00719_));
 sky130_fd_sc_hd__inv_2 _13557_ (.A(\CPU_Xreg_value_a4[9][0] ),
    .Y(_07733_));
 sky130_fd_sc_hd__nor2_4 _13558_ (.A(_07733_),
    .B(_07654_),
    .Y(_07734_));
 sky130_fd_sc_hd__a211o_4 _13559_ (.A1(_07188_),
    .A2(_07654_),
    .B1(_07530_),
    .C1(_07734_),
    .X(_00718_));
 sky130_fd_sc_hd__or2_4 _13560_ (.A(_06986_),
    .B(_07537_),
    .X(_07735_));
 sky130_fd_sc_hd__nor2_4 _13561_ (.A(_07449_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__buf_2 _13562_ (.A(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__buf_2 _13563_ (.A(_07737_),
    .X(_07738_));
 sky130_fd_sc_hd__buf_2 _13564_ (.A(_07702_),
    .X(_07739_));
 sky130_fd_sc_hd__buf_2 _13565_ (.A(_07737_),
    .X(_07740_));
 sky130_fd_sc_hd__nor2_4 _13566_ (.A(\CPU_Xreg_value_a4[10][31] ),
    .B(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__a211o_4 _13567_ (.A1(_07535_),
    .A2(_07738_),
    .B1(_07739_),
    .C1(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__inv_2 _13568_ (.A(_07742_),
    .Y(_00717_));
 sky130_fd_sc_hd__nor2_4 _13569_ (.A(\CPU_Xreg_value_a4[10][30] ),
    .B(_07740_),
    .Y(_07743_));
 sky130_fd_sc_hd__a211o_4 _13570_ (.A1(_07545_),
    .A2(_07738_),
    .B1(_07739_),
    .C1(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__inv_2 _13571_ (.A(_07744_),
    .Y(_00716_));
 sky130_fd_sc_hd__buf_2 _13572_ (.A(_07736_),
    .X(_07745_));
 sky130_fd_sc_hd__buf_2 _13573_ (.A(_07745_),
    .X(_07746_));
 sky130_fd_sc_hd__buf_2 _13574_ (.A(_07737_),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_4 _13575_ (.A(\CPU_Xreg_value_a4[10][29] ),
    .B(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__a211o_4 _13576_ (.A1(_07549_),
    .A2(_07746_),
    .B1(_07739_),
    .C1(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__inv_2 _13577_ (.A(_07749_),
    .Y(_00715_));
 sky130_fd_sc_hd__nor2_4 _13578_ (.A(\CPU_Xreg_value_a4[10][28] ),
    .B(_07747_),
    .Y(_07750_));
 sky130_fd_sc_hd__a211o_4 _13579_ (.A1(_07552_),
    .A2(_07746_),
    .B1(_07739_),
    .C1(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__inv_2 _13580_ (.A(_07751_),
    .Y(_00714_));
 sky130_fd_sc_hd__nor2_4 _13581_ (.A(\CPU_Xreg_value_a4[10][27] ),
    .B(_07747_),
    .Y(_07752_));
 sky130_fd_sc_hd__a211o_4 _13582_ (.A1(_07556_),
    .A2(_07746_),
    .B1(_07739_),
    .C1(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__inv_2 _13583_ (.A(_07753_),
    .Y(_00713_));
 sky130_fd_sc_hd__nor2_4 _13584_ (.A(\CPU_Xreg_value_a4[10][26] ),
    .B(_07747_),
    .Y(_07754_));
 sky130_fd_sc_hd__a211o_4 _13585_ (.A1(_07561_),
    .A2(_07746_),
    .B1(_07739_),
    .C1(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__inv_2 _13586_ (.A(_07755_),
    .Y(_00712_));
 sky130_fd_sc_hd__buf_2 _13587_ (.A(_07702_),
    .X(_07756_));
 sky130_fd_sc_hd__nor2_4 _13588_ (.A(\CPU_Xreg_value_a4[10][25] ),
    .B(_07747_),
    .Y(_07757_));
 sky130_fd_sc_hd__a211o_4 _13589_ (.A1(_07564_),
    .A2(_07746_),
    .B1(_07756_),
    .C1(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__inv_2 _13590_ (.A(_07758_),
    .Y(_00711_));
 sky130_fd_sc_hd__nor2_4 _13591_ (.A(\CPU_Xreg_value_a4[10][24] ),
    .B(_07747_),
    .Y(_07759_));
 sky130_fd_sc_hd__a211o_4 _13592_ (.A1(_07567_),
    .A2(_07746_),
    .B1(_07756_),
    .C1(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__inv_2 _13593_ (.A(_07760_),
    .Y(_00710_));
 sky130_fd_sc_hd__buf_2 _13594_ (.A(_07745_),
    .X(_07761_));
 sky130_fd_sc_hd__buf_2 _13595_ (.A(_07737_),
    .X(_07762_));
 sky130_fd_sc_hd__nor2_4 _13596_ (.A(\CPU_Xreg_value_a4[10][23] ),
    .B(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__a211o_4 _13597_ (.A1(_07571_),
    .A2(_07761_),
    .B1(_07756_),
    .C1(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__inv_2 _13598_ (.A(_07764_),
    .Y(_00709_));
 sky130_fd_sc_hd__nor2_4 _13599_ (.A(\CPU_Xreg_value_a4[10][22] ),
    .B(_07762_),
    .Y(_07765_));
 sky130_fd_sc_hd__a211o_4 _13600_ (.A1(_07574_),
    .A2(_07761_),
    .B1(_07756_),
    .C1(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__inv_2 _13601_ (.A(_07766_),
    .Y(_00708_));
 sky130_fd_sc_hd__nor2_4 _13602_ (.A(\CPU_Xreg_value_a4[10][21] ),
    .B(_07762_),
    .Y(_07767_));
 sky130_fd_sc_hd__a211o_4 _13603_ (.A1(_07578_),
    .A2(_07761_),
    .B1(_07756_),
    .C1(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__inv_2 _13604_ (.A(_07768_),
    .Y(_00707_));
 sky130_fd_sc_hd__nor2_4 _13605_ (.A(\CPU_Xreg_value_a4[10][20] ),
    .B(_07762_),
    .Y(_07769_));
 sky130_fd_sc_hd__a211o_4 _13606_ (.A1(_07582_),
    .A2(_07761_),
    .B1(_07756_),
    .C1(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__inv_2 _13607_ (.A(_07770_),
    .Y(_00706_));
 sky130_fd_sc_hd__buf_2 _13608_ (.A(_07702_),
    .X(_07771_));
 sky130_fd_sc_hd__nor2_4 _13609_ (.A(\CPU_Xreg_value_a4[10][19] ),
    .B(_07762_),
    .Y(_07772_));
 sky130_fd_sc_hd__a211o_4 _13610_ (.A1(_07585_),
    .A2(_07761_),
    .B1(_07771_),
    .C1(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__inv_2 _13611_ (.A(_07773_),
    .Y(_00705_));
 sky130_fd_sc_hd__nor2_4 _13612_ (.A(\CPU_Xreg_value_a4[10][18] ),
    .B(_07762_),
    .Y(_07774_));
 sky130_fd_sc_hd__a211o_4 _13613_ (.A1(_07588_),
    .A2(_07761_),
    .B1(_07771_),
    .C1(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__inv_2 _13614_ (.A(_07775_),
    .Y(_00704_));
 sky130_fd_sc_hd__buf_2 _13615_ (.A(_07737_),
    .X(_07776_));
 sky130_fd_sc_hd__buf_2 _13616_ (.A(_07736_),
    .X(_07777_));
 sky130_fd_sc_hd__nor2_4 _13617_ (.A(\CPU_Xreg_value_a4[10][17] ),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__a211o_4 _13618_ (.A1(_07593_),
    .A2(_07776_),
    .B1(_07771_),
    .C1(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__inv_2 _13619_ (.A(_07779_),
    .Y(_00703_));
 sky130_fd_sc_hd__nor2_4 _13620_ (.A(\CPU_Xreg_value_a4[10][16] ),
    .B(_07777_),
    .Y(_07780_));
 sky130_fd_sc_hd__a211o_4 _13621_ (.A1(_07596_),
    .A2(_07776_),
    .B1(_07771_),
    .C1(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__inv_2 _13622_ (.A(_07781_),
    .Y(_00702_));
 sky130_fd_sc_hd__nor2_4 _13623_ (.A(\CPU_Xreg_value_a4[10][15] ),
    .B(_07777_),
    .Y(_07782_));
 sky130_fd_sc_hd__a211o_4 _13624_ (.A1(_07600_),
    .A2(_07776_),
    .B1(_07771_),
    .C1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__inv_2 _13625_ (.A(_07783_),
    .Y(_00701_));
 sky130_fd_sc_hd__nor2_4 _13626_ (.A(\CPU_Xreg_value_a4[10][14] ),
    .B(_07777_),
    .Y(_07784_));
 sky130_fd_sc_hd__a211o_4 _13627_ (.A1(_07604_),
    .A2(_07776_),
    .B1(_07771_),
    .C1(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__inv_2 _13628_ (.A(_07785_),
    .Y(_00700_));
 sky130_fd_sc_hd__buf_2 _13629_ (.A(_07702_),
    .X(_07786_));
 sky130_fd_sc_hd__nor2_4 _13630_ (.A(\CPU_Xreg_value_a4[10][13] ),
    .B(_07777_),
    .Y(_07787_));
 sky130_fd_sc_hd__a211o_4 _13631_ (.A1(_07607_),
    .A2(_07776_),
    .B1(_07786_),
    .C1(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__inv_2 _13632_ (.A(_07788_),
    .Y(_00699_));
 sky130_fd_sc_hd__nor2_4 _13633_ (.A(\CPU_Xreg_value_a4[10][12] ),
    .B(_07777_),
    .Y(_07789_));
 sky130_fd_sc_hd__a211o_4 _13634_ (.A1(_07610_),
    .A2(_07776_),
    .B1(_07786_),
    .C1(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__inv_2 _13635_ (.A(_07790_),
    .Y(_00698_));
 sky130_fd_sc_hd__buf_2 _13636_ (.A(_07737_),
    .X(_07791_));
 sky130_fd_sc_hd__buf_2 _13637_ (.A(_07736_),
    .X(_07792_));
 sky130_fd_sc_hd__nor2_4 _13638_ (.A(\CPU_Xreg_value_a4[10][11] ),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__a211o_4 _13639_ (.A1(_07614_),
    .A2(_07791_),
    .B1(_07786_),
    .C1(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__inv_2 _13640_ (.A(_07794_),
    .Y(_00697_));
 sky130_fd_sc_hd__nor2_4 _13641_ (.A(\CPU_Xreg_value_a4[10][10] ),
    .B(_07792_),
    .Y(_07795_));
 sky130_fd_sc_hd__a211o_4 _13642_ (.A1(_07617_),
    .A2(_07791_),
    .B1(_07786_),
    .C1(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__inv_2 _13643_ (.A(_07796_),
    .Y(_00696_));
 sky130_fd_sc_hd__nor2_4 _13644_ (.A(\CPU_Xreg_value_a4[10][9] ),
    .B(_07792_),
    .Y(_07797_));
 sky130_fd_sc_hd__a211o_4 _13645_ (.A1(_07621_),
    .A2(_07791_),
    .B1(_07786_),
    .C1(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__inv_2 _13646_ (.A(_07798_),
    .Y(_00695_));
 sky130_fd_sc_hd__nor2_4 _13647_ (.A(\CPU_Xreg_value_a4[10][8] ),
    .B(_07792_),
    .Y(_07799_));
 sky130_fd_sc_hd__a211o_4 _13648_ (.A1(_07625_),
    .A2(_07791_),
    .B1(_07786_),
    .C1(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__inv_2 _13649_ (.A(_07800_),
    .Y(_00694_));
 sky130_fd_sc_hd__buf_2 _13650_ (.A(CPU_reset_a3),
    .X(_07801_));
 sky130_fd_sc_hd__buf_2 _13651_ (.A(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__buf_2 _13652_ (.A(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__nor2_4 _13653_ (.A(\CPU_Xreg_value_a4[10][7] ),
    .B(_07792_),
    .Y(_07804_));
 sky130_fd_sc_hd__a211o_4 _13654_ (.A1(_07628_),
    .A2(_07791_),
    .B1(_07803_),
    .C1(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__inv_2 _13655_ (.A(_07805_),
    .Y(_00693_));
 sky130_fd_sc_hd__nor2_4 _13656_ (.A(\CPU_Xreg_value_a4[10][6] ),
    .B(_07792_),
    .Y(_07806_));
 sky130_fd_sc_hd__a211o_4 _13657_ (.A1(_07631_),
    .A2(_07791_),
    .B1(_07803_),
    .C1(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__inv_2 _13658_ (.A(_07807_),
    .Y(_00692_));
 sky130_fd_sc_hd__nor2_4 _13659_ (.A(\CPU_Xreg_value_a4[10][5] ),
    .B(_07745_),
    .Y(_07808_));
 sky130_fd_sc_hd__a211o_4 _13660_ (.A1(_07635_),
    .A2(_07740_),
    .B1(_07803_),
    .C1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__inv_2 _13661_ (.A(_07809_),
    .Y(_00691_));
 sky130_fd_sc_hd__nor2_4 _13662_ (.A(\CPU_Xreg_value_a4[10][4] ),
    .B(_07745_),
    .Y(_07810_));
 sky130_fd_sc_hd__a211o_4 _13663_ (.A1(_07638_),
    .A2(_07740_),
    .B1(_07803_),
    .C1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__inv_2 _13664_ (.A(_07811_),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _13665_ (.A(\CPU_Xreg_value_a4[10][3] ),
    .Y(_07812_));
 sky130_fd_sc_hd__nor2_4 _13666_ (.A(_07812_),
    .B(_07738_),
    .Y(_07813_));
 sky130_fd_sc_hd__a211o_4 _13667_ (.A1(_07642_),
    .A2(_07738_),
    .B1(_07530_),
    .C1(_07813_),
    .X(_00689_));
 sky130_fd_sc_hd__nor2_4 _13668_ (.A(\CPU_Xreg_value_a4[10][2] ),
    .B(_07745_),
    .Y(_07814_));
 sky130_fd_sc_hd__a211o_4 _13669_ (.A1(_07093_),
    .A2(_07740_),
    .B1(_07803_),
    .C1(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__inv_2 _13670_ (.A(_07815_),
    .Y(_00688_));
 sky130_fd_sc_hd__buf_2 _13671_ (.A(_07273_),
    .X(_07816_));
 sky130_fd_sc_hd__inv_2 _13672_ (.A(\CPU_Xreg_value_a4[10][1] ),
    .Y(_07817_));
 sky130_fd_sc_hd__nor2_4 _13673_ (.A(_07817_),
    .B(_07738_),
    .Y(_07818_));
 sky130_fd_sc_hd__a211o_4 _13674_ (.A1(_07097_),
    .A2(_07738_),
    .B1(_07816_),
    .C1(_07818_),
    .X(_00687_));
 sky130_fd_sc_hd__nor2_4 _13675_ (.A(\CPU_Xreg_value_a4[10][0] ),
    .B(_07745_),
    .Y(_07819_));
 sky130_fd_sc_hd__a211o_4 _13676_ (.A1(_07101_),
    .A2(_07740_),
    .B1(_07803_),
    .C1(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__inv_2 _13677_ (.A(_07820_),
    .Y(_00686_));
 sky130_fd_sc_hd__or2_4 _13678_ (.A(_07104_),
    .B(_07537_),
    .X(_07821_));
 sky130_fd_sc_hd__nor2_4 _13679_ (.A(_07449_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__buf_2 _13680_ (.A(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__buf_2 _13681_ (.A(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__buf_2 _13682_ (.A(_07802_),
    .X(_07825_));
 sky130_fd_sc_hd__buf_2 _13683_ (.A(_07822_),
    .X(_07826_));
 sky130_fd_sc_hd__buf_2 _13684_ (.A(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__nor2_4 _13685_ (.A(\CPU_Xreg_value_a4[11][31] ),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__a211o_4 _13686_ (.A1(_07535_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__inv_2 _13687_ (.A(_07829_),
    .Y(_00685_));
 sky130_fd_sc_hd__buf_2 _13688_ (.A(_07826_),
    .X(_07830_));
 sky130_fd_sc_hd__nor2_4 _13689_ (.A(\CPU_Xreg_value_a4[11][30] ),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__a211o_4 _13690_ (.A1(_07545_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__inv_2 _13691_ (.A(_07832_),
    .Y(_00684_));
 sky130_fd_sc_hd__nor2_4 _13692_ (.A(\CPU_Xreg_value_a4[11][29] ),
    .B(_07830_),
    .Y(_07833_));
 sky130_fd_sc_hd__a211o_4 _13693_ (.A1(_07549_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__inv_2 _13694_ (.A(_07834_),
    .Y(_00683_));
 sky130_fd_sc_hd__nor2_4 _13695_ (.A(\CPU_Xreg_value_a4[11][28] ),
    .B(_07830_),
    .Y(_07835_));
 sky130_fd_sc_hd__a211o_4 _13696_ (.A1(_07552_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__inv_2 _13697_ (.A(_07836_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_4 _13698_ (.A(\CPU_Xreg_value_a4[11][27] ),
    .B(_07830_),
    .Y(_07837_));
 sky130_fd_sc_hd__a211o_4 _13699_ (.A1(_07556_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07837_),
    .X(_07838_));
 sky130_fd_sc_hd__inv_2 _13700_ (.A(_07838_),
    .Y(_00681_));
 sky130_fd_sc_hd__nor2_4 _13701_ (.A(\CPU_Xreg_value_a4[11][26] ),
    .B(_07830_),
    .Y(_07839_));
 sky130_fd_sc_hd__a211o_4 _13702_ (.A1(_07561_),
    .A2(_07824_),
    .B1(_07825_),
    .C1(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__inv_2 _13703_ (.A(_07840_),
    .Y(_00680_));
 sky130_fd_sc_hd__buf_2 _13704_ (.A(_07826_),
    .X(_07841_));
 sky130_fd_sc_hd__buf_2 _13705_ (.A(_07802_),
    .X(_07842_));
 sky130_fd_sc_hd__nor2_4 _13706_ (.A(\CPU_Xreg_value_a4[11][25] ),
    .B(_07830_),
    .Y(_07843_));
 sky130_fd_sc_hd__a211o_4 _13707_ (.A1(_07564_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__inv_2 _13708_ (.A(_07844_),
    .Y(_00679_));
 sky130_fd_sc_hd__buf_2 _13709_ (.A(_07826_),
    .X(_07845_));
 sky130_fd_sc_hd__nor2_4 _13710_ (.A(\CPU_Xreg_value_a4[11][24] ),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__a211o_4 _13711_ (.A1(_07567_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__inv_2 _13712_ (.A(_07847_),
    .Y(_00678_));
 sky130_fd_sc_hd__nor2_4 _13713_ (.A(\CPU_Xreg_value_a4[11][23] ),
    .B(_07845_),
    .Y(_07848_));
 sky130_fd_sc_hd__a211o_4 _13714_ (.A1(_07571_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__inv_2 _13715_ (.A(_07849_),
    .Y(_00677_));
 sky130_fd_sc_hd__nor2_4 _13716_ (.A(\CPU_Xreg_value_a4[11][22] ),
    .B(_07845_),
    .Y(_07850_));
 sky130_fd_sc_hd__a211o_4 _13717_ (.A1(_07574_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__inv_2 _13718_ (.A(_07851_),
    .Y(_00676_));
 sky130_fd_sc_hd__nor2_4 _13719_ (.A(\CPU_Xreg_value_a4[11][21] ),
    .B(_07845_),
    .Y(_07852_));
 sky130_fd_sc_hd__a211o_4 _13720_ (.A1(_07578_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__inv_2 _13721_ (.A(_07853_),
    .Y(_00675_));
 sky130_fd_sc_hd__nor2_4 _13722_ (.A(\CPU_Xreg_value_a4[11][20] ),
    .B(_07845_),
    .Y(_07854_));
 sky130_fd_sc_hd__a211o_4 _13723_ (.A1(_07582_),
    .A2(_07841_),
    .B1(_07842_),
    .C1(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__inv_2 _13724_ (.A(_07855_),
    .Y(_00674_));
 sky130_fd_sc_hd__buf_2 _13725_ (.A(_07826_),
    .X(_07856_));
 sky130_fd_sc_hd__buf_2 _13726_ (.A(_07802_),
    .X(_07857_));
 sky130_fd_sc_hd__nor2_4 _13727_ (.A(\CPU_Xreg_value_a4[11][19] ),
    .B(_07845_),
    .Y(_07858_));
 sky130_fd_sc_hd__a211o_4 _13728_ (.A1(_07585_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__inv_2 _13729_ (.A(_07859_),
    .Y(_00673_));
 sky130_fd_sc_hd__buf_2 _13730_ (.A(_07822_),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_4 _13731_ (.A(\CPU_Xreg_value_a4[11][18] ),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__a211o_4 _13732_ (.A1(_07588_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__inv_2 _13733_ (.A(_07862_),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_4 _13734_ (.A(\CPU_Xreg_value_a4[11][17] ),
    .B(_07860_),
    .Y(_07863_));
 sky130_fd_sc_hd__a211o_4 _13735_ (.A1(_07593_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__inv_2 _13736_ (.A(_07864_),
    .Y(_00671_));
 sky130_fd_sc_hd__nor2_4 _13737_ (.A(\CPU_Xreg_value_a4[11][16] ),
    .B(_07860_),
    .Y(_07865_));
 sky130_fd_sc_hd__a211o_4 _13738_ (.A1(_07596_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__inv_2 _13739_ (.A(_07866_),
    .Y(_00670_));
 sky130_fd_sc_hd__nor2_4 _13740_ (.A(\CPU_Xreg_value_a4[11][15] ),
    .B(_07860_),
    .Y(_07867_));
 sky130_fd_sc_hd__a211o_4 _13741_ (.A1(_07600_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__inv_2 _13742_ (.A(_07868_),
    .Y(_00669_));
 sky130_fd_sc_hd__nor2_4 _13743_ (.A(\CPU_Xreg_value_a4[11][14] ),
    .B(_07860_),
    .Y(_07869_));
 sky130_fd_sc_hd__a211o_4 _13744_ (.A1(_07604_),
    .A2(_07856_),
    .B1(_07857_),
    .C1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__inv_2 _13745_ (.A(_07870_),
    .Y(_00668_));
 sky130_fd_sc_hd__buf_2 _13746_ (.A(_07826_),
    .X(_07871_));
 sky130_fd_sc_hd__buf_2 _13747_ (.A(_07802_),
    .X(_07872_));
 sky130_fd_sc_hd__nor2_4 _13748_ (.A(\CPU_Xreg_value_a4[11][13] ),
    .B(_07860_),
    .Y(_07873_));
 sky130_fd_sc_hd__a211o_4 _13749_ (.A1(_07607_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__inv_2 _13750_ (.A(_07874_),
    .Y(_00667_));
 sky130_fd_sc_hd__buf_2 _13751_ (.A(_07822_),
    .X(_07875_));
 sky130_fd_sc_hd__nor2_4 _13752_ (.A(\CPU_Xreg_value_a4[11][12] ),
    .B(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__a211o_4 _13753_ (.A1(_07610_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__inv_2 _13754_ (.A(_07877_),
    .Y(_00666_));
 sky130_fd_sc_hd__nor2_4 _13755_ (.A(\CPU_Xreg_value_a4[11][11] ),
    .B(_07875_),
    .Y(_07878_));
 sky130_fd_sc_hd__a211o_4 _13756_ (.A1(_07614_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__inv_2 _13757_ (.A(_07879_),
    .Y(_00665_));
 sky130_fd_sc_hd__nor2_4 _13758_ (.A(\CPU_Xreg_value_a4[11][10] ),
    .B(_07875_),
    .Y(_07880_));
 sky130_fd_sc_hd__a211o_4 _13759_ (.A1(_07617_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__inv_2 _13760_ (.A(_07881_),
    .Y(_00664_));
 sky130_fd_sc_hd__nor2_4 _13761_ (.A(\CPU_Xreg_value_a4[11][9] ),
    .B(_07875_),
    .Y(_07882_));
 sky130_fd_sc_hd__a211o_4 _13762_ (.A1(_07621_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__inv_2 _13763_ (.A(_07883_),
    .Y(_00663_));
 sky130_fd_sc_hd__nor2_4 _13764_ (.A(\CPU_Xreg_value_a4[11][8] ),
    .B(_07875_),
    .Y(_07884_));
 sky130_fd_sc_hd__a211o_4 _13765_ (.A1(_07625_),
    .A2(_07871_),
    .B1(_07872_),
    .C1(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__inv_2 _13766_ (.A(_07885_),
    .Y(_00662_));
 sky130_fd_sc_hd__buf_2 _13767_ (.A(_07802_),
    .X(_07886_));
 sky130_fd_sc_hd__nor2_4 _13768_ (.A(\CPU_Xreg_value_a4[11][7] ),
    .B(_07875_),
    .Y(_07887_));
 sky130_fd_sc_hd__a211o_4 _13769_ (.A1(_07628_),
    .A2(_07827_),
    .B1(_07886_),
    .C1(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__inv_2 _13770_ (.A(_07888_),
    .Y(_00661_));
 sky130_fd_sc_hd__nor2_4 _13771_ (.A(\CPU_Xreg_value_a4[11][6] ),
    .B(_07823_),
    .Y(_07889_));
 sky130_fd_sc_hd__a211o_4 _13772_ (.A1(_07631_),
    .A2(_07827_),
    .B1(_07886_),
    .C1(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__inv_2 _13773_ (.A(_07890_),
    .Y(_00660_));
 sky130_fd_sc_hd__nor2_4 _13774_ (.A(\CPU_Xreg_value_a4[11][5] ),
    .B(_07823_),
    .Y(_07891_));
 sky130_fd_sc_hd__a211o_4 _13775_ (.A1(_07635_),
    .A2(_07827_),
    .B1(_07886_),
    .C1(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__inv_2 _13776_ (.A(_07892_),
    .Y(_00659_));
 sky130_fd_sc_hd__nor2_4 _13777_ (.A(\CPU_Xreg_value_a4[11][4] ),
    .B(_07823_),
    .Y(_07893_));
 sky130_fd_sc_hd__a211o_4 _13778_ (.A1(_07638_),
    .A2(_07827_),
    .B1(_07886_),
    .C1(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__inv_2 _13779_ (.A(_07894_),
    .Y(_00658_));
 sky130_fd_sc_hd__buf_2 _13780_ (.A(_07823_),
    .X(_07895_));
 sky130_fd_sc_hd__inv_2 _13781_ (.A(\CPU_Xreg_value_a4[11][3] ),
    .Y(_07896_));
 sky130_fd_sc_hd__nor2_4 _13782_ (.A(_07896_),
    .B(_07895_),
    .Y(_07897_));
 sky130_fd_sc_hd__a211o_4 _13783_ (.A1(_07642_),
    .A2(_07895_),
    .B1(_07816_),
    .C1(_07897_),
    .X(_00657_));
 sky130_fd_sc_hd__nor2_4 _13784_ (.A(\CPU_Xreg_value_a4[11][2] ),
    .B(_07823_),
    .Y(_07898_));
 sky130_fd_sc_hd__a211o_4 _13785_ (.A1(_07093_),
    .A2(_07827_),
    .B1(_07886_),
    .C1(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__inv_2 _13786_ (.A(_07899_),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_2 _13787_ (.A(\CPU_Xreg_value_a4[11][1] ),
    .Y(_07900_));
 sky130_fd_sc_hd__nor2_4 _13788_ (.A(_07900_),
    .B(_07895_),
    .Y(_07901_));
 sky130_fd_sc_hd__a211o_4 _13789_ (.A1(_07097_),
    .A2(_07895_),
    .B1(_07816_),
    .C1(_07901_),
    .X(_00655_));
 sky130_fd_sc_hd__inv_2 _13790_ (.A(\CPU_Xreg_value_a4[11][0] ),
    .Y(_07902_));
 sky130_fd_sc_hd__nor2_4 _13791_ (.A(_07902_),
    .B(_07895_),
    .Y(_07903_));
 sky130_fd_sc_hd__a211o_4 _13792_ (.A1(_07188_),
    .A2(_07895_),
    .B1(_07816_),
    .C1(_07903_),
    .X(_00654_));
 sky130_fd_sc_hd__or2_4 _13793_ (.A(_07191_),
    .B(_07536_),
    .X(_07904_));
 sky130_fd_sc_hd__or2_4 _13794_ (.A(_06156_),
    .B(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__nor2_4 _13795_ (.A(_07449_),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__buf_2 _13796_ (.A(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__buf_2 _13797_ (.A(_07907_),
    .X(_07908_));
 sky130_fd_sc_hd__buf_2 _13798_ (.A(_07907_),
    .X(_07909_));
 sky130_fd_sc_hd__nor2_4 _13799_ (.A(\CPU_Xreg_value_a4[12][31] ),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__a211o_4 _13800_ (.A1(_07535_),
    .A2(_07908_),
    .B1(_07886_),
    .C1(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__inv_2 _13801_ (.A(_07911_),
    .Y(_00653_));
 sky130_fd_sc_hd__buf_2 _13802_ (.A(_07801_),
    .X(_07912_));
 sky130_fd_sc_hd__buf_2 _13803_ (.A(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__nor2_4 _13804_ (.A(\CPU_Xreg_value_a4[12][30] ),
    .B(_07909_),
    .Y(_07914_));
 sky130_fd_sc_hd__a211o_4 _13805_ (.A1(_07545_),
    .A2(_07908_),
    .B1(_07913_),
    .C1(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__inv_2 _13806_ (.A(_07915_),
    .Y(_00652_));
 sky130_fd_sc_hd__buf_2 _13807_ (.A(_07906_),
    .X(_07916_));
 sky130_fd_sc_hd__buf_2 _13808_ (.A(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__buf_2 _13809_ (.A(_07907_),
    .X(_07918_));
 sky130_fd_sc_hd__nor2_4 _13810_ (.A(\CPU_Xreg_value_a4[12][29] ),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__a211o_4 _13811_ (.A1(_07549_),
    .A2(_07917_),
    .B1(_07913_),
    .C1(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__inv_2 _13812_ (.A(_07920_),
    .Y(_00651_));
 sky130_fd_sc_hd__nor2_4 _13813_ (.A(\CPU_Xreg_value_a4[12][28] ),
    .B(_07918_),
    .Y(_07921_));
 sky130_fd_sc_hd__a211o_4 _13814_ (.A1(_07552_),
    .A2(_07917_),
    .B1(_07913_),
    .C1(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__inv_2 _13815_ (.A(_07922_),
    .Y(_00650_));
 sky130_fd_sc_hd__nor2_4 _13816_ (.A(\CPU_Xreg_value_a4[12][27] ),
    .B(_07918_),
    .Y(_07923_));
 sky130_fd_sc_hd__a211o_4 _13817_ (.A1(_07556_),
    .A2(_07917_),
    .B1(_07913_),
    .C1(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__inv_2 _13818_ (.A(_07924_),
    .Y(_00649_));
 sky130_fd_sc_hd__nor2_4 _13819_ (.A(\CPU_Xreg_value_a4[12][26] ),
    .B(_07918_),
    .Y(_07925_));
 sky130_fd_sc_hd__a211o_4 _13820_ (.A1(_07561_),
    .A2(_07917_),
    .B1(_07913_),
    .C1(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__inv_2 _13821_ (.A(_07926_),
    .Y(_00648_));
 sky130_fd_sc_hd__nor2_4 _13822_ (.A(\CPU_Xreg_value_a4[12][25] ),
    .B(_07918_),
    .Y(_07927_));
 sky130_fd_sc_hd__a211o_4 _13823_ (.A1(_07564_),
    .A2(_07917_),
    .B1(_07913_),
    .C1(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__inv_2 _13824_ (.A(_07928_),
    .Y(_00647_));
 sky130_fd_sc_hd__buf_2 _13825_ (.A(_07912_),
    .X(_07929_));
 sky130_fd_sc_hd__nor2_4 _13826_ (.A(\CPU_Xreg_value_a4[12][24] ),
    .B(_07918_),
    .Y(_07930_));
 sky130_fd_sc_hd__a211o_4 _13827_ (.A1(_07567_),
    .A2(_07917_),
    .B1(_07929_),
    .C1(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__inv_2 _13828_ (.A(_07931_),
    .Y(_00646_));
 sky130_fd_sc_hd__buf_2 _13829_ (.A(_07916_),
    .X(_07932_));
 sky130_fd_sc_hd__buf_2 _13830_ (.A(_07907_),
    .X(_07933_));
 sky130_fd_sc_hd__nor2_4 _13831_ (.A(\CPU_Xreg_value_a4[12][23] ),
    .B(_07933_),
    .Y(_07934_));
 sky130_fd_sc_hd__a211o_4 _13832_ (.A1(_07571_),
    .A2(_07932_),
    .B1(_07929_),
    .C1(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__inv_2 _13833_ (.A(_07935_),
    .Y(_00645_));
 sky130_fd_sc_hd__nor2_4 _13834_ (.A(\CPU_Xreg_value_a4[12][22] ),
    .B(_07933_),
    .Y(_07936_));
 sky130_fd_sc_hd__a211o_4 _13835_ (.A1(_07574_),
    .A2(_07932_),
    .B1(_07929_),
    .C1(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__inv_2 _13836_ (.A(_07937_),
    .Y(_00644_));
 sky130_fd_sc_hd__nor2_4 _13837_ (.A(\CPU_Xreg_value_a4[12][21] ),
    .B(_07933_),
    .Y(_07938_));
 sky130_fd_sc_hd__a211o_4 _13838_ (.A1(_07578_),
    .A2(_07932_),
    .B1(_07929_),
    .C1(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__inv_2 _13839_ (.A(_07939_),
    .Y(_00643_));
 sky130_fd_sc_hd__nor2_4 _13840_ (.A(\CPU_Xreg_value_a4[12][20] ),
    .B(_07933_),
    .Y(_07940_));
 sky130_fd_sc_hd__a211o_4 _13841_ (.A1(_07582_),
    .A2(_07932_),
    .B1(_07929_),
    .C1(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__inv_2 _13842_ (.A(_07941_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor2_4 _13843_ (.A(\CPU_Xreg_value_a4[12][19] ),
    .B(_07933_),
    .Y(_07942_));
 sky130_fd_sc_hd__a211o_4 _13844_ (.A1(_07585_),
    .A2(_07932_),
    .B1(_07929_),
    .C1(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__inv_2 _13845_ (.A(_07943_),
    .Y(_00641_));
 sky130_fd_sc_hd__buf_2 _13846_ (.A(_07912_),
    .X(_07944_));
 sky130_fd_sc_hd__nor2_4 _13847_ (.A(\CPU_Xreg_value_a4[12][18] ),
    .B(_07933_),
    .Y(_07945_));
 sky130_fd_sc_hd__a211o_4 _13848_ (.A1(_07588_),
    .A2(_07932_),
    .B1(_07944_),
    .C1(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__inv_2 _13849_ (.A(_07946_),
    .Y(_00640_));
 sky130_fd_sc_hd__buf_2 _13850_ (.A(_07907_),
    .X(_07947_));
 sky130_fd_sc_hd__buf_2 _13851_ (.A(_07906_),
    .X(_07948_));
 sky130_fd_sc_hd__nor2_4 _13852_ (.A(\CPU_Xreg_value_a4[12][17] ),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__a211o_4 _13853_ (.A1(_07593_),
    .A2(_07947_),
    .B1(_07944_),
    .C1(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__inv_2 _13854_ (.A(_07950_),
    .Y(_00639_));
 sky130_fd_sc_hd__nor2_4 _13855_ (.A(\CPU_Xreg_value_a4[12][16] ),
    .B(_07948_),
    .Y(_07951_));
 sky130_fd_sc_hd__a211o_4 _13856_ (.A1(_07596_),
    .A2(_07947_),
    .B1(_07944_),
    .C1(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__inv_2 _13857_ (.A(_07952_),
    .Y(_00638_));
 sky130_fd_sc_hd__nor2_4 _13858_ (.A(\CPU_Xreg_value_a4[12][15] ),
    .B(_07948_),
    .Y(_07953_));
 sky130_fd_sc_hd__a211o_4 _13859_ (.A1(_07600_),
    .A2(_07947_),
    .B1(_07944_),
    .C1(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__inv_2 _13860_ (.A(_07954_),
    .Y(_00637_));
 sky130_fd_sc_hd__nor2_4 _13861_ (.A(\CPU_Xreg_value_a4[12][14] ),
    .B(_07948_),
    .Y(_07955_));
 sky130_fd_sc_hd__a211o_4 _13862_ (.A1(_07604_),
    .A2(_07947_),
    .B1(_07944_),
    .C1(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__inv_2 _13863_ (.A(_07956_),
    .Y(_00636_));
 sky130_fd_sc_hd__nor2_4 _13864_ (.A(\CPU_Xreg_value_a4[12][13] ),
    .B(_07948_),
    .Y(_07957_));
 sky130_fd_sc_hd__a211o_4 _13865_ (.A1(_07607_),
    .A2(_07947_),
    .B1(_07944_),
    .C1(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__inv_2 _13866_ (.A(_07958_),
    .Y(_00635_));
 sky130_fd_sc_hd__buf_2 _13867_ (.A(_07912_),
    .X(_07959_));
 sky130_fd_sc_hd__nor2_4 _13868_ (.A(\CPU_Xreg_value_a4[12][12] ),
    .B(_07948_),
    .Y(_07960_));
 sky130_fd_sc_hd__a211o_4 _13869_ (.A1(_07610_),
    .A2(_07947_),
    .B1(_07959_),
    .C1(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__inv_2 _13870_ (.A(_07961_),
    .Y(_00634_));
 sky130_fd_sc_hd__buf_2 _13871_ (.A(_07907_),
    .X(_07962_));
 sky130_fd_sc_hd__buf_2 _13872_ (.A(_07906_),
    .X(_07963_));
 sky130_fd_sc_hd__nor2_4 _13873_ (.A(\CPU_Xreg_value_a4[12][11] ),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__a211o_4 _13874_ (.A1(_07614_),
    .A2(_07962_),
    .B1(_07959_),
    .C1(_07964_),
    .X(_07965_));
 sky130_fd_sc_hd__inv_2 _13875_ (.A(_07965_),
    .Y(_00633_));
 sky130_fd_sc_hd__nor2_4 _13876_ (.A(\CPU_Xreg_value_a4[12][10] ),
    .B(_07963_),
    .Y(_07966_));
 sky130_fd_sc_hd__a211o_4 _13877_ (.A1(_07617_),
    .A2(_07962_),
    .B1(_07959_),
    .C1(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__inv_2 _13878_ (.A(_07967_),
    .Y(_00632_));
 sky130_fd_sc_hd__nor2_4 _13879_ (.A(\CPU_Xreg_value_a4[12][9] ),
    .B(_07963_),
    .Y(_07968_));
 sky130_fd_sc_hd__a211o_4 _13880_ (.A1(_07621_),
    .A2(_07962_),
    .B1(_07959_),
    .C1(_07968_),
    .X(_07969_));
 sky130_fd_sc_hd__inv_2 _13881_ (.A(_07969_),
    .Y(_00631_));
 sky130_fd_sc_hd__nor2_4 _13882_ (.A(\CPU_Xreg_value_a4[12][8] ),
    .B(_07963_),
    .Y(_07970_));
 sky130_fd_sc_hd__a211o_4 _13883_ (.A1(_07625_),
    .A2(_07962_),
    .B1(_07959_),
    .C1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__inv_2 _13884_ (.A(_07971_),
    .Y(_00630_));
 sky130_fd_sc_hd__nor2_4 _13885_ (.A(\CPU_Xreg_value_a4[12][7] ),
    .B(_07963_),
    .Y(_07972_));
 sky130_fd_sc_hd__a211o_4 _13886_ (.A1(_07628_),
    .A2(_07962_),
    .B1(_07959_),
    .C1(_07972_),
    .X(_07973_));
 sky130_fd_sc_hd__inv_2 _13887_ (.A(_07973_),
    .Y(_00629_));
 sky130_fd_sc_hd__buf_2 _13888_ (.A(_07912_),
    .X(_07974_));
 sky130_fd_sc_hd__nor2_4 _13889_ (.A(\CPU_Xreg_value_a4[12][6] ),
    .B(_07963_),
    .Y(_07975_));
 sky130_fd_sc_hd__a211o_4 _13890_ (.A1(_07631_),
    .A2(_07962_),
    .B1(_07974_),
    .C1(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__inv_2 _13891_ (.A(_07976_),
    .Y(_00628_));
 sky130_fd_sc_hd__nor2_4 _13892_ (.A(\CPU_Xreg_value_a4[12][5] ),
    .B(_07916_),
    .Y(_07977_));
 sky130_fd_sc_hd__a211o_4 _13893_ (.A1(_07635_),
    .A2(_07909_),
    .B1(_07974_),
    .C1(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__inv_2 _13894_ (.A(_07978_),
    .Y(_00627_));
 sky130_fd_sc_hd__nor2_4 _13895_ (.A(\CPU_Xreg_value_a4[12][4] ),
    .B(_07916_),
    .Y(_07979_));
 sky130_fd_sc_hd__a211o_4 _13896_ (.A1(_07638_),
    .A2(_07909_),
    .B1(_07974_),
    .C1(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__inv_2 _13897_ (.A(_07980_),
    .Y(_00626_));
 sky130_fd_sc_hd__inv_2 _13898_ (.A(\CPU_Xreg_value_a4[12][3] ),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_4 _13899_ (.A(_07981_),
    .B(_07908_),
    .Y(_07982_));
 sky130_fd_sc_hd__a211o_4 _13900_ (.A1(_07642_),
    .A2(_07908_),
    .B1(_07816_),
    .C1(_07982_),
    .X(_00625_));
 sky130_fd_sc_hd__inv_2 _13901_ (.A(\CPU_Xreg_value_a4[12][2] ),
    .Y(_07983_));
 sky130_fd_sc_hd__nor2_4 _13902_ (.A(_07983_),
    .B(_07908_),
    .Y(_07984_));
 sky130_fd_sc_hd__a211o_4 _13903_ (.A1(_07272_),
    .A2(_07908_),
    .B1(_07816_),
    .C1(_07984_),
    .X(_00624_));
 sky130_fd_sc_hd__nor2_4 _13904_ (.A(\CPU_Xreg_value_a4[12][1] ),
    .B(_07916_),
    .Y(_07985_));
 sky130_fd_sc_hd__a211o_4 _13905_ (.A1(_07277_),
    .A2(_07909_),
    .B1(_07974_),
    .C1(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__inv_2 _13906_ (.A(_07986_),
    .Y(_00623_));
 sky130_fd_sc_hd__nor2_4 _13907_ (.A(\CPU_Xreg_value_a4[12][0] ),
    .B(_07916_),
    .Y(_07987_));
 sky130_fd_sc_hd__a211o_4 _13908_ (.A1(_07101_),
    .A2(_07909_),
    .B1(_07974_),
    .C1(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__inv_2 _13909_ (.A(_07988_),
    .Y(_00622_));
 sky130_fd_sc_hd__or2_4 _13910_ (.A(_06152_),
    .B(_07904_),
    .X(_07989_));
 sky130_fd_sc_hd__or2_4 _13911_ (.A(_06165_),
    .B(_07989_),
    .X(_07990_));
 sky130_fd_sc_hd__inv_2 _13912_ (.A(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__buf_2 _13913_ (.A(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__buf_2 _13914_ (.A(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__buf_2 _13915_ (.A(_07991_),
    .X(_07994_));
 sky130_fd_sc_hd__nor2_4 _13916_ (.A(\CPU_Xreg_value_a4[13][31] ),
    .B(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__a211o_4 _13917_ (.A1(_07535_),
    .A2(_07993_),
    .B1(_07974_),
    .C1(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__inv_2 _13918_ (.A(_07996_),
    .Y(_00621_));
 sky130_fd_sc_hd__buf_2 _13919_ (.A(_07912_),
    .X(_07997_));
 sky130_fd_sc_hd__nor2_4 _13920_ (.A(\CPU_Xreg_value_a4[13][30] ),
    .B(_07994_),
    .Y(_07998_));
 sky130_fd_sc_hd__a211o_4 _13921_ (.A1(_07545_),
    .A2(_07993_),
    .B1(_07997_),
    .C1(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__inv_2 _13922_ (.A(_07999_),
    .Y(_00620_));
 sky130_fd_sc_hd__nor2_4 _13923_ (.A(\CPU_Xreg_value_a4[13][29] ),
    .B(_07994_),
    .Y(_08000_));
 sky130_fd_sc_hd__a211o_4 _13924_ (.A1(_07549_),
    .A2(_07993_),
    .B1(_07997_),
    .C1(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__inv_2 _13925_ (.A(_08001_),
    .Y(_00619_));
 sky130_fd_sc_hd__buf_2 _13926_ (.A(_07992_),
    .X(_08002_));
 sky130_fd_sc_hd__nor2_4 _13927_ (.A(\CPU_Xreg_value_a4[13][28] ),
    .B(_07994_),
    .Y(_08003_));
 sky130_fd_sc_hd__a211o_4 _13928_ (.A1(_07552_),
    .A2(_08002_),
    .B1(_07997_),
    .C1(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__inv_2 _13929_ (.A(_08004_),
    .Y(_00618_));
 sky130_fd_sc_hd__buf_2 _13930_ (.A(_07991_),
    .X(_08005_));
 sky130_fd_sc_hd__nor2_4 _13931_ (.A(\CPU_Xreg_value_a4[13][27] ),
    .B(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__a211o_4 _13932_ (.A1(_07556_),
    .A2(_08002_),
    .B1(_07997_),
    .C1(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__inv_2 _13933_ (.A(_08007_),
    .Y(_00617_));
 sky130_fd_sc_hd__nor2_4 _13934_ (.A(\CPU_Xreg_value_a4[13][26] ),
    .B(_08005_),
    .Y(_08008_));
 sky130_fd_sc_hd__a211o_4 _13935_ (.A1(_07561_),
    .A2(_08002_),
    .B1(_07997_),
    .C1(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__inv_2 _13936_ (.A(_08009_),
    .Y(_00616_));
 sky130_fd_sc_hd__nor2_4 _13937_ (.A(\CPU_Xreg_value_a4[13][25] ),
    .B(_08005_),
    .Y(_08010_));
 sky130_fd_sc_hd__a211o_4 _13938_ (.A1(_07564_),
    .A2(_08002_),
    .B1(_07997_),
    .C1(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__inv_2 _13939_ (.A(_08011_),
    .Y(_00615_));
 sky130_fd_sc_hd__buf_2 _13940_ (.A(_07801_),
    .X(_08012_));
 sky130_fd_sc_hd__buf_2 _13941_ (.A(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__nor2_4 _13942_ (.A(\CPU_Xreg_value_a4[13][24] ),
    .B(_08005_),
    .Y(_08014_));
 sky130_fd_sc_hd__a211o_4 _13943_ (.A1(_07567_),
    .A2(_08002_),
    .B1(_08013_),
    .C1(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__inv_2 _13944_ (.A(_08015_),
    .Y(_00614_));
 sky130_fd_sc_hd__nor2_4 _13945_ (.A(\CPU_Xreg_value_a4[13][23] ),
    .B(_08005_),
    .Y(_08016_));
 sky130_fd_sc_hd__a211o_4 _13946_ (.A1(_07571_),
    .A2(_08002_),
    .B1(_08013_),
    .C1(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__inv_2 _13947_ (.A(_08017_),
    .Y(_00613_));
 sky130_fd_sc_hd__buf_2 _13948_ (.A(_07992_),
    .X(_08018_));
 sky130_fd_sc_hd__nor2_4 _13949_ (.A(\CPU_Xreg_value_a4[13][22] ),
    .B(_08005_),
    .Y(_08019_));
 sky130_fd_sc_hd__a211o_4 _13950_ (.A1(_07574_),
    .A2(_08018_),
    .B1(_08013_),
    .C1(_08019_),
    .X(_08020_));
 sky130_fd_sc_hd__inv_2 _13951_ (.A(_08020_),
    .Y(_00612_));
 sky130_fd_sc_hd__buf_2 _13952_ (.A(_07991_),
    .X(_08021_));
 sky130_fd_sc_hd__nor2_4 _13953_ (.A(\CPU_Xreg_value_a4[13][21] ),
    .B(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__a211o_4 _13954_ (.A1(_07578_),
    .A2(_08018_),
    .B1(_08013_),
    .C1(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__inv_2 _13955_ (.A(_08023_),
    .Y(_00611_));
 sky130_fd_sc_hd__nor2_4 _13956_ (.A(\CPU_Xreg_value_a4[13][20] ),
    .B(_08021_),
    .Y(_08024_));
 sky130_fd_sc_hd__a211o_4 _13957_ (.A1(_07582_),
    .A2(_08018_),
    .B1(_08013_),
    .C1(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__inv_2 _13958_ (.A(_08025_),
    .Y(_00610_));
 sky130_fd_sc_hd__nor2_4 _13959_ (.A(\CPU_Xreg_value_a4[13][19] ),
    .B(_08021_),
    .Y(_08026_));
 sky130_fd_sc_hd__a211o_4 _13960_ (.A1(_07585_),
    .A2(_08018_),
    .B1(_08013_),
    .C1(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__inv_2 _13961_ (.A(_08027_),
    .Y(_00609_));
 sky130_fd_sc_hd__buf_2 _13962_ (.A(_08012_),
    .X(_08028_));
 sky130_fd_sc_hd__nor2_4 _13963_ (.A(\CPU_Xreg_value_a4[13][18] ),
    .B(_08021_),
    .Y(_08029_));
 sky130_fd_sc_hd__a211o_4 _13964_ (.A1(_07588_),
    .A2(_08018_),
    .B1(_08028_),
    .C1(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__inv_2 _13965_ (.A(_08030_),
    .Y(_00608_));
 sky130_fd_sc_hd__nor2_4 _13966_ (.A(\CPU_Xreg_value_a4[13][17] ),
    .B(_08021_),
    .Y(_08031_));
 sky130_fd_sc_hd__a211o_4 _13967_ (.A1(_07593_),
    .A2(_08018_),
    .B1(_08028_),
    .C1(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__inv_2 _13968_ (.A(_08032_),
    .Y(_00607_));
 sky130_fd_sc_hd__buf_2 _13969_ (.A(_07992_),
    .X(_08033_));
 sky130_fd_sc_hd__nor2_4 _13970_ (.A(\CPU_Xreg_value_a4[13][16] ),
    .B(_08021_),
    .Y(_08034_));
 sky130_fd_sc_hd__a211o_4 _13971_ (.A1(_07596_),
    .A2(_08033_),
    .B1(_08028_),
    .C1(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__inv_2 _13972_ (.A(_08035_),
    .Y(_00606_));
 sky130_fd_sc_hd__buf_2 _13973_ (.A(_07991_),
    .X(_08036_));
 sky130_fd_sc_hd__nor2_4 _13974_ (.A(\CPU_Xreg_value_a4[13][15] ),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__a211o_4 _13975_ (.A1(_07600_),
    .A2(_08033_),
    .B1(_08028_),
    .C1(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__inv_2 _13976_ (.A(_08038_),
    .Y(_00605_));
 sky130_fd_sc_hd__nor2_4 _13977_ (.A(\CPU_Xreg_value_a4[13][14] ),
    .B(_08036_),
    .Y(_08039_));
 sky130_fd_sc_hd__a211o_4 _13978_ (.A1(_07604_),
    .A2(_08033_),
    .B1(_08028_),
    .C1(_08039_),
    .X(_08040_));
 sky130_fd_sc_hd__inv_2 _13979_ (.A(_08040_),
    .Y(_00604_));
 sky130_fd_sc_hd__nor2_4 _13980_ (.A(\CPU_Xreg_value_a4[13][13] ),
    .B(_08036_),
    .Y(_08041_));
 sky130_fd_sc_hd__a211o_4 _13981_ (.A1(_07607_),
    .A2(_08033_),
    .B1(_08028_),
    .C1(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__inv_2 _13982_ (.A(_08042_),
    .Y(_00603_));
 sky130_fd_sc_hd__buf_2 _13983_ (.A(_08012_),
    .X(_08043_));
 sky130_fd_sc_hd__nor2_4 _13984_ (.A(\CPU_Xreg_value_a4[13][12] ),
    .B(_08036_),
    .Y(_08044_));
 sky130_fd_sc_hd__a211o_4 _13985_ (.A1(_07610_),
    .A2(_08033_),
    .B1(_08043_),
    .C1(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__inv_2 _13986_ (.A(_08045_),
    .Y(_00602_));
 sky130_fd_sc_hd__nor2_4 _13987_ (.A(\CPU_Xreg_value_a4[13][11] ),
    .B(_08036_),
    .Y(_08046_));
 sky130_fd_sc_hd__a211o_4 _13988_ (.A1(_07614_),
    .A2(_08033_),
    .B1(_08043_),
    .C1(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__inv_2 _13989_ (.A(_08047_),
    .Y(_00601_));
 sky130_fd_sc_hd__buf_2 _13990_ (.A(_07992_),
    .X(_08048_));
 sky130_fd_sc_hd__nor2_4 _13991_ (.A(\CPU_Xreg_value_a4[13][10] ),
    .B(_08036_),
    .Y(_08049_));
 sky130_fd_sc_hd__a211o_4 _13992_ (.A1(_07617_),
    .A2(_08048_),
    .B1(_08043_),
    .C1(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__inv_2 _13993_ (.A(_08050_),
    .Y(_00600_));
 sky130_fd_sc_hd__buf_2 _13994_ (.A(_07991_),
    .X(_08051_));
 sky130_fd_sc_hd__nor2_4 _13995_ (.A(\CPU_Xreg_value_a4[13][9] ),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__a211o_4 _13996_ (.A1(_07621_),
    .A2(_08048_),
    .B1(_08043_),
    .C1(_08052_),
    .X(_08053_));
 sky130_fd_sc_hd__inv_2 _13997_ (.A(_08053_),
    .Y(_00599_));
 sky130_fd_sc_hd__nor2_4 _13998_ (.A(\CPU_Xreg_value_a4[13][8] ),
    .B(_08051_),
    .Y(_08054_));
 sky130_fd_sc_hd__a211o_4 _13999_ (.A1(_07625_),
    .A2(_08048_),
    .B1(_08043_),
    .C1(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__inv_2 _14000_ (.A(_08055_),
    .Y(_00598_));
 sky130_fd_sc_hd__nor2_4 _14001_ (.A(\CPU_Xreg_value_a4[13][7] ),
    .B(_08051_),
    .Y(_08056_));
 sky130_fd_sc_hd__a211o_4 _14002_ (.A1(_07628_),
    .A2(_08048_),
    .B1(_08043_),
    .C1(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__inv_2 _14003_ (.A(_08057_),
    .Y(_00597_));
 sky130_fd_sc_hd__buf_2 _14004_ (.A(_08012_),
    .X(_08058_));
 sky130_fd_sc_hd__nor2_4 _14005_ (.A(\CPU_Xreg_value_a4[13][6] ),
    .B(_08051_),
    .Y(_08059_));
 sky130_fd_sc_hd__a211o_4 _14006_ (.A1(_07631_),
    .A2(_08048_),
    .B1(_08058_),
    .C1(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__inv_2 _14007_ (.A(_08060_),
    .Y(_00596_));
 sky130_fd_sc_hd__nor2_4 _14008_ (.A(\CPU_Xreg_value_a4[13][5] ),
    .B(_08051_),
    .Y(_08061_));
 sky130_fd_sc_hd__a211o_4 _14009_ (.A1(_07635_),
    .A2(_08048_),
    .B1(_08058_),
    .C1(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__inv_2 _14010_ (.A(_08062_),
    .Y(_00595_));
 sky130_fd_sc_hd__nor2_4 _14011_ (.A(\CPU_Xreg_value_a4[13][4] ),
    .B(_08051_),
    .Y(_08063_));
 sky130_fd_sc_hd__a211o_4 _14012_ (.A1(_07638_),
    .A2(_07994_),
    .B1(_08058_),
    .C1(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__inv_2 _14013_ (.A(_08064_),
    .Y(_00594_));
 sky130_fd_sc_hd__buf_2 _14014_ (.A(_06101_),
    .X(_08065_));
 sky130_fd_sc_hd__buf_2 _14015_ (.A(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__and2_4 _14016_ (.A(\CPU_Xreg_value_a4[13][3] ),
    .B(_07990_),
    .X(_08067_));
 sky130_fd_sc_hd__a211o_4 _14017_ (.A1(_07642_),
    .A2(_07993_),
    .B1(_08066_),
    .C1(_08067_),
    .X(_00593_));
 sky130_fd_sc_hd__and2_4 _14018_ (.A(\CPU_Xreg_value_a4[13][2] ),
    .B(_07990_),
    .X(_08068_));
 sky130_fd_sc_hd__a211o_4 _14019_ (.A1(_07272_),
    .A2(_07993_),
    .B1(_08066_),
    .C1(_08068_),
    .X(_00592_));
 sky130_fd_sc_hd__nor2_4 _14020_ (.A(\CPU_Xreg_value_a4[13][1] ),
    .B(_07992_),
    .Y(_08069_));
 sky130_fd_sc_hd__a211o_4 _14021_ (.A1(_07277_),
    .A2(_07994_),
    .B1(_08058_),
    .C1(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__inv_2 _14022_ (.A(_08070_),
    .Y(_00591_));
 sky130_fd_sc_hd__and2_4 _14023_ (.A(\CPU_Xreg_value_a4[13][0] ),
    .B(_07990_),
    .X(_08071_));
 sky130_fd_sc_hd__a211o_4 _14024_ (.A1(_07188_),
    .A2(_07993_),
    .B1(_08066_),
    .C1(_08071_),
    .X(_00590_));
 sky130_fd_sc_hd__buf_2 _14025_ (.A(_06503_),
    .X(_08072_));
 sky130_fd_sc_hd__or2_4 _14026_ (.A(_06986_),
    .B(_07904_),
    .X(_08073_));
 sky130_fd_sc_hd__nor2_4 _14027_ (.A(_06165_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__buf_2 _14028_ (.A(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__buf_2 _14029_ (.A(_08075_),
    .X(_08076_));
 sky130_fd_sc_hd__buf_2 _14030_ (.A(_08074_),
    .X(_08077_));
 sky130_fd_sc_hd__buf_2 _14031_ (.A(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__nor2_4 _14032_ (.A(\CPU_Xreg_value_a4[14][31] ),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__a211o_4 _14033_ (.A1(_08072_),
    .A2(_08076_),
    .B1(_08058_),
    .C1(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__inv_2 _14034_ (.A(_08080_),
    .Y(_00589_));
 sky130_fd_sc_hd__buf_2 _14035_ (.A(_06515_),
    .X(_08081_));
 sky130_fd_sc_hd__buf_2 _14036_ (.A(_08077_),
    .X(_08082_));
 sky130_fd_sc_hd__nor2_4 _14037_ (.A(\CPU_Xreg_value_a4[14][30] ),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__a211o_4 _14038_ (.A1(_08081_),
    .A2(_08076_),
    .B1(_08058_),
    .C1(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__inv_2 _14039_ (.A(_08084_),
    .Y(_00588_));
 sky130_fd_sc_hd__buf_2 _14040_ (.A(_06531_),
    .X(_08085_));
 sky130_fd_sc_hd__buf_2 _14041_ (.A(_08012_),
    .X(_08086_));
 sky130_fd_sc_hd__nor2_4 _14042_ (.A(\CPU_Xreg_value_a4[14][29] ),
    .B(_08082_),
    .Y(_08087_));
 sky130_fd_sc_hd__a211o_4 _14043_ (.A1(_08085_),
    .A2(_08076_),
    .B1(_08086_),
    .C1(_08087_),
    .X(_08088_));
 sky130_fd_sc_hd__inv_2 _14044_ (.A(_08088_),
    .Y(_00587_));
 sky130_fd_sc_hd__buf_2 _14045_ (.A(_06539_),
    .X(_08089_));
 sky130_fd_sc_hd__nor2_4 _14046_ (.A(\CPU_Xreg_value_a4[14][28] ),
    .B(_08082_),
    .Y(_08090_));
 sky130_fd_sc_hd__a211o_4 _14047_ (.A1(_08089_),
    .A2(_08076_),
    .B1(_08086_),
    .C1(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__inv_2 _14048_ (.A(_08091_),
    .Y(_00586_));
 sky130_fd_sc_hd__buf_2 _14049_ (.A(_06564_),
    .X(_08092_));
 sky130_fd_sc_hd__nor2_4 _14050_ (.A(\CPU_Xreg_value_a4[14][27] ),
    .B(_08082_),
    .Y(_08093_));
 sky130_fd_sc_hd__a211o_4 _14051_ (.A1(_08092_),
    .A2(_08076_),
    .B1(_08086_),
    .C1(_08093_),
    .X(_08094_));
 sky130_fd_sc_hd__inv_2 _14052_ (.A(_08094_),
    .Y(_00585_));
 sky130_fd_sc_hd__buf_2 _14053_ (.A(_06574_),
    .X(_08095_));
 sky130_fd_sc_hd__nor2_4 _14054_ (.A(\CPU_Xreg_value_a4[14][26] ),
    .B(_08082_),
    .Y(_08096_));
 sky130_fd_sc_hd__a211o_4 _14055_ (.A1(_08095_),
    .A2(_08076_),
    .B1(_08086_),
    .C1(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__inv_2 _14056_ (.A(_08097_),
    .Y(_00584_));
 sky130_fd_sc_hd__buf_2 _14057_ (.A(_06589_),
    .X(_08098_));
 sky130_fd_sc_hd__buf_2 _14058_ (.A(_08077_),
    .X(_08099_));
 sky130_fd_sc_hd__nor2_4 _14059_ (.A(\CPU_Xreg_value_a4[14][25] ),
    .B(_08082_),
    .Y(_08100_));
 sky130_fd_sc_hd__a211o_4 _14060_ (.A1(_08098_),
    .A2(_08099_),
    .B1(_08086_),
    .C1(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__inv_2 _14061_ (.A(_08101_),
    .Y(_00583_));
 sky130_fd_sc_hd__buf_2 _14062_ (.A(_06599_),
    .X(_08102_));
 sky130_fd_sc_hd__buf_2 _14063_ (.A(_08077_),
    .X(_08103_));
 sky130_fd_sc_hd__nor2_4 _14064_ (.A(\CPU_Xreg_value_a4[14][24] ),
    .B(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__a211o_4 _14065_ (.A1(_08102_),
    .A2(_08099_),
    .B1(_08086_),
    .C1(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__inv_2 _14066_ (.A(_08105_),
    .Y(_00582_));
 sky130_fd_sc_hd__buf_2 _14067_ (.A(_06619_),
    .X(_08106_));
 sky130_fd_sc_hd__buf_2 _14068_ (.A(_08012_),
    .X(_08107_));
 sky130_fd_sc_hd__nor2_4 _14069_ (.A(\CPU_Xreg_value_a4[14][23] ),
    .B(_08103_),
    .Y(_08108_));
 sky130_fd_sc_hd__a211o_4 _14070_ (.A1(_08106_),
    .A2(_08099_),
    .B1(_08107_),
    .C1(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__inv_2 _14071_ (.A(_08109_),
    .Y(_00581_));
 sky130_fd_sc_hd__buf_2 _14072_ (.A(_06627_),
    .X(_08110_));
 sky130_fd_sc_hd__nor2_4 _14073_ (.A(\CPU_Xreg_value_a4[14][22] ),
    .B(_08103_),
    .Y(_08111_));
 sky130_fd_sc_hd__a211o_4 _14074_ (.A1(_08110_),
    .A2(_08099_),
    .B1(_08107_),
    .C1(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__inv_2 _14075_ (.A(_08112_),
    .Y(_00580_));
 sky130_fd_sc_hd__buf_2 _14076_ (.A(_06642_),
    .X(_08113_));
 sky130_fd_sc_hd__nor2_4 _14077_ (.A(\CPU_Xreg_value_a4[14][21] ),
    .B(_08103_),
    .Y(_08114_));
 sky130_fd_sc_hd__a211o_4 _14078_ (.A1(_08113_),
    .A2(_08099_),
    .B1(_08107_),
    .C1(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__inv_2 _14079_ (.A(_08115_),
    .Y(_00579_));
 sky130_fd_sc_hd__buf_2 _14080_ (.A(_06651_),
    .X(_08116_));
 sky130_fd_sc_hd__nor2_4 _14081_ (.A(\CPU_Xreg_value_a4[14][20] ),
    .B(_08103_),
    .Y(_08117_));
 sky130_fd_sc_hd__a211o_4 _14082_ (.A1(_08116_),
    .A2(_08099_),
    .B1(_08107_),
    .C1(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__inv_2 _14083_ (.A(_08118_),
    .Y(_00578_));
 sky130_fd_sc_hd__buf_2 _14084_ (.A(_06673_),
    .X(_08119_));
 sky130_fd_sc_hd__buf_2 _14085_ (.A(_08077_),
    .X(_08120_));
 sky130_fd_sc_hd__nor2_4 _14086_ (.A(\CPU_Xreg_value_a4[14][19] ),
    .B(_08103_),
    .Y(_08121_));
 sky130_fd_sc_hd__a211o_4 _14087_ (.A1(_08119_),
    .A2(_08120_),
    .B1(_08107_),
    .C1(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__inv_2 _14088_ (.A(_08122_),
    .Y(_00577_));
 sky130_fd_sc_hd__buf_2 _14089_ (.A(_06682_),
    .X(_08123_));
 sky130_fd_sc_hd__buf_2 _14090_ (.A(_08074_),
    .X(_08124_));
 sky130_fd_sc_hd__nor2_4 _14091_ (.A(\CPU_Xreg_value_a4[14][18] ),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__a211o_4 _14092_ (.A1(_08123_),
    .A2(_08120_),
    .B1(_08107_),
    .C1(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__inv_2 _14093_ (.A(_08126_),
    .Y(_00576_));
 sky130_fd_sc_hd__buf_2 _14094_ (.A(_06692_),
    .X(_08127_));
 sky130_fd_sc_hd__buf_2 _14095_ (.A(_07801_),
    .X(_08128_));
 sky130_fd_sc_hd__buf_2 _14096_ (.A(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__nor2_4 _14097_ (.A(\CPU_Xreg_value_a4[14][17] ),
    .B(_08124_),
    .Y(_08130_));
 sky130_fd_sc_hd__a211o_4 _14098_ (.A1(_08127_),
    .A2(_08120_),
    .B1(_08129_),
    .C1(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__inv_2 _14099_ (.A(_08131_),
    .Y(_00575_));
 sky130_fd_sc_hd__buf_2 _14100_ (.A(_06701_),
    .X(_08132_));
 sky130_fd_sc_hd__nor2_4 _14101_ (.A(\CPU_Xreg_value_a4[14][16] ),
    .B(_08124_),
    .Y(_08133_));
 sky130_fd_sc_hd__a211o_4 _14102_ (.A1(_08132_),
    .A2(_08120_),
    .B1(_08129_),
    .C1(_08133_),
    .X(_08134_));
 sky130_fd_sc_hd__inv_2 _14103_ (.A(_08134_),
    .Y(_00574_));
 sky130_fd_sc_hd__buf_2 _14104_ (.A(_06724_),
    .X(_08135_));
 sky130_fd_sc_hd__nor2_4 _14105_ (.A(\CPU_Xreg_value_a4[14][15] ),
    .B(_08124_),
    .Y(_08136_));
 sky130_fd_sc_hd__a211o_4 _14106_ (.A1(_08135_),
    .A2(_08120_),
    .B1(_08129_),
    .C1(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__inv_2 _14107_ (.A(_08137_),
    .Y(_00573_));
 sky130_fd_sc_hd__buf_2 _14108_ (.A(_06733_),
    .X(_08138_));
 sky130_fd_sc_hd__nor2_4 _14109_ (.A(\CPU_Xreg_value_a4[14][14] ),
    .B(_08124_),
    .Y(_08139_));
 sky130_fd_sc_hd__a211o_4 _14110_ (.A1(_08138_),
    .A2(_08120_),
    .B1(_08129_),
    .C1(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__inv_2 _14111_ (.A(_08140_),
    .Y(_00572_));
 sky130_fd_sc_hd__buf_2 _14112_ (.A(_06743_),
    .X(_08141_));
 sky130_fd_sc_hd__buf_2 _14113_ (.A(_08077_),
    .X(_08142_));
 sky130_fd_sc_hd__nor2_4 _14114_ (.A(\CPU_Xreg_value_a4[14][13] ),
    .B(_08124_),
    .Y(_08143_));
 sky130_fd_sc_hd__a211o_4 _14115_ (.A1(_08141_),
    .A2(_08142_),
    .B1(_08129_),
    .C1(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__inv_2 _14116_ (.A(_08144_),
    .Y(_00571_));
 sky130_fd_sc_hd__buf_2 _14117_ (.A(_06752_),
    .X(_08145_));
 sky130_fd_sc_hd__buf_2 _14118_ (.A(_08074_),
    .X(_08146_));
 sky130_fd_sc_hd__nor2_4 _14119_ (.A(\CPU_Xreg_value_a4[14][12] ),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__a211o_4 _14120_ (.A1(_08145_),
    .A2(_08142_),
    .B1(_08129_),
    .C1(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__inv_2 _14121_ (.A(_08148_),
    .Y(_00570_));
 sky130_fd_sc_hd__buf_2 _14122_ (.A(_06770_),
    .X(_08149_));
 sky130_fd_sc_hd__buf_2 _14123_ (.A(_08128_),
    .X(_08150_));
 sky130_fd_sc_hd__nor2_4 _14124_ (.A(\CPU_Xreg_value_a4[14][11] ),
    .B(_08146_),
    .Y(_08151_));
 sky130_fd_sc_hd__a211o_4 _14125_ (.A1(_08149_),
    .A2(_08142_),
    .B1(_08150_),
    .C1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__inv_2 _14126_ (.A(_08152_),
    .Y(_00569_));
 sky130_fd_sc_hd__buf_2 _14127_ (.A(_06778_),
    .X(_08153_));
 sky130_fd_sc_hd__nor2_4 _14128_ (.A(\CPU_Xreg_value_a4[14][10] ),
    .B(_08146_),
    .Y(_08154_));
 sky130_fd_sc_hd__a211o_4 _14129_ (.A1(_08153_),
    .A2(_08142_),
    .B1(_08150_),
    .C1(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__inv_2 _14130_ (.A(_08155_),
    .Y(_00568_));
 sky130_fd_sc_hd__buf_2 _14131_ (.A(_06791_),
    .X(_08156_));
 sky130_fd_sc_hd__nor2_4 _14132_ (.A(\CPU_Xreg_value_a4[14][9] ),
    .B(_08146_),
    .Y(_08157_));
 sky130_fd_sc_hd__a211o_4 _14133_ (.A1(_08156_),
    .A2(_08142_),
    .B1(_08150_),
    .C1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__inv_2 _14134_ (.A(_08158_),
    .Y(_00567_));
 sky130_fd_sc_hd__buf_2 _14135_ (.A(_06799_),
    .X(_08159_));
 sky130_fd_sc_hd__nor2_4 _14136_ (.A(\CPU_Xreg_value_a4[14][8] ),
    .B(_08146_),
    .Y(_08160_));
 sky130_fd_sc_hd__a211o_4 _14137_ (.A1(_08159_),
    .A2(_08142_),
    .B1(_08150_),
    .C1(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__inv_2 _14138_ (.A(_08161_),
    .Y(_00566_));
 sky130_fd_sc_hd__buf_2 _14139_ (.A(_06820_),
    .X(_08162_));
 sky130_fd_sc_hd__nor2_4 _14140_ (.A(\CPU_Xreg_value_a4[14][7] ),
    .B(_08146_),
    .Y(_08163_));
 sky130_fd_sc_hd__a211o_4 _14141_ (.A1(_08162_),
    .A2(_08078_),
    .B1(_08150_),
    .C1(_08163_),
    .X(_08164_));
 sky130_fd_sc_hd__inv_2 _14142_ (.A(_08164_),
    .Y(_00565_));
 sky130_fd_sc_hd__buf_2 _14143_ (.A(_06828_),
    .X(_08165_));
 sky130_fd_sc_hd__nor2_4 _14144_ (.A(\CPU_Xreg_value_a4[14][6] ),
    .B(_08075_),
    .Y(_08166_));
 sky130_fd_sc_hd__a211o_4 _14145_ (.A1(_08165_),
    .A2(_08078_),
    .B1(_08150_),
    .C1(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__inv_2 _14146_ (.A(_08167_),
    .Y(_00564_));
 sky130_fd_sc_hd__buf_2 _14147_ (.A(_06837_),
    .X(_08168_));
 sky130_fd_sc_hd__buf_2 _14148_ (.A(_08128_),
    .X(_08169_));
 sky130_fd_sc_hd__nor2_4 _14149_ (.A(\CPU_Xreg_value_a4[14][5] ),
    .B(_08075_),
    .Y(_08170_));
 sky130_fd_sc_hd__a211o_4 _14150_ (.A1(_08168_),
    .A2(_08078_),
    .B1(_08169_),
    .C1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__inv_2 _14151_ (.A(_08171_),
    .Y(_00563_));
 sky130_fd_sc_hd__nor2_4 _14152_ (.A(\CPU_Xreg_value_a4[14][4] ),
    .B(_08075_),
    .Y(_08172_));
 sky130_fd_sc_hd__a211o_4 _14153_ (.A1(_06843_),
    .A2(_08078_),
    .B1(_08169_),
    .C1(_08172_),
    .X(_08173_));
 sky130_fd_sc_hd__inv_2 _14154_ (.A(_08173_),
    .Y(_00562_));
 sky130_fd_sc_hd__buf_2 _14155_ (.A(_07641_),
    .X(_08174_));
 sky130_fd_sc_hd__buf_2 _14156_ (.A(_08075_),
    .X(_08175_));
 sky130_fd_sc_hd__inv_2 _14157_ (.A(\CPU_Xreg_value_a4[14][3] ),
    .Y(_08176_));
 sky130_fd_sc_hd__nor2_4 _14158_ (.A(_08176_),
    .B(_08175_),
    .Y(_08177_));
 sky130_fd_sc_hd__a211o_4 _14159_ (.A1(_08174_),
    .A2(_08175_),
    .B1(_08066_),
    .C1(_08177_),
    .X(_00561_));
 sky130_fd_sc_hd__buf_2 _14160_ (.A(_07271_),
    .X(_08178_));
 sky130_fd_sc_hd__inv_2 _14161_ (.A(\CPU_Xreg_value_a4[14][2] ),
    .Y(_08179_));
 sky130_fd_sc_hd__nor2_4 _14162_ (.A(_08179_),
    .B(_08175_),
    .Y(_08180_));
 sky130_fd_sc_hd__a211o_4 _14163_ (.A1(_08178_),
    .A2(_08175_),
    .B1(_08066_),
    .C1(_08180_),
    .X(_00560_));
 sky130_fd_sc_hd__buf_2 _14164_ (.A(_07096_),
    .X(_08181_));
 sky130_fd_sc_hd__inv_2 _14165_ (.A(\CPU_Xreg_value_a4[14][1] ),
    .Y(_08182_));
 sky130_fd_sc_hd__nor2_4 _14166_ (.A(_08182_),
    .B(_08175_),
    .Y(_08183_));
 sky130_fd_sc_hd__a211o_4 _14167_ (.A1(_08181_),
    .A2(_08175_),
    .B1(_08066_),
    .C1(_08183_),
    .X(_00559_));
 sky130_fd_sc_hd__buf_2 _14168_ (.A(_07100_),
    .X(_08184_));
 sky130_fd_sc_hd__nor2_4 _14169_ (.A(\CPU_Xreg_value_a4[14][0] ),
    .B(_08075_),
    .Y(_08185_));
 sky130_fd_sc_hd__a211o_4 _14170_ (.A1(_08184_),
    .A2(_08078_),
    .B1(_08169_),
    .C1(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__inv_2 _14171_ (.A(_08186_),
    .Y(_00558_));
 sky130_fd_sc_hd__or2_4 _14172_ (.A(_07104_),
    .B(_07904_),
    .X(_08187_));
 sky130_fd_sc_hd__nor2_4 _14173_ (.A(_06165_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__buf_2 _14174_ (.A(_08188_),
    .X(_08189_));
 sky130_fd_sc_hd__buf_2 _14175_ (.A(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__buf_2 _14176_ (.A(_08189_),
    .X(_08191_));
 sky130_fd_sc_hd__nor2_4 _14177_ (.A(\CPU_Xreg_value_a4[15][31] ),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__a211o_4 _14178_ (.A1(_08072_),
    .A2(_08190_),
    .B1(_08169_),
    .C1(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__inv_2 _14179_ (.A(_08193_),
    .Y(_00557_));
 sky130_fd_sc_hd__nor2_4 _14180_ (.A(\CPU_Xreg_value_a4[15][30] ),
    .B(_08191_),
    .Y(_08194_));
 sky130_fd_sc_hd__a211o_4 _14181_ (.A1(_08081_),
    .A2(_08190_),
    .B1(_08169_),
    .C1(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__inv_2 _14182_ (.A(_08195_),
    .Y(_00556_));
 sky130_fd_sc_hd__nor2_4 _14183_ (.A(\CPU_Xreg_value_a4[15][29] ),
    .B(_08191_),
    .Y(_08196_));
 sky130_fd_sc_hd__a211o_4 _14184_ (.A1(_08085_),
    .A2(_08190_),
    .B1(_08169_),
    .C1(_08196_),
    .X(_08197_));
 sky130_fd_sc_hd__inv_2 _14185_ (.A(_08197_),
    .Y(_00555_));
 sky130_fd_sc_hd__buf_2 _14186_ (.A(_08128_),
    .X(_08198_));
 sky130_fd_sc_hd__nor2_4 _14187_ (.A(\CPU_Xreg_value_a4[15][28] ),
    .B(_08191_),
    .Y(_08199_));
 sky130_fd_sc_hd__a211o_4 _14188_ (.A1(_08089_),
    .A2(_08190_),
    .B1(_08198_),
    .C1(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__inv_2 _14189_ (.A(_08200_),
    .Y(_00554_));
 sky130_fd_sc_hd__buf_2 _14190_ (.A(_08188_),
    .X(_08201_));
 sky130_fd_sc_hd__buf_2 _14191_ (.A(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__nor2_4 _14192_ (.A(\CPU_Xreg_value_a4[15][27] ),
    .B(_08191_),
    .Y(_08203_));
 sky130_fd_sc_hd__a211o_4 _14193_ (.A1(_08092_),
    .A2(_08202_),
    .B1(_08198_),
    .C1(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__inv_2 _14194_ (.A(_08204_),
    .Y(_00553_));
 sky130_fd_sc_hd__nor2_4 _14195_ (.A(\CPU_Xreg_value_a4[15][26] ),
    .B(_08191_),
    .Y(_08205_));
 sky130_fd_sc_hd__a211o_4 _14196_ (.A1(_08095_),
    .A2(_08202_),
    .B1(_08198_),
    .C1(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__inv_2 _14197_ (.A(_08206_),
    .Y(_00552_));
 sky130_fd_sc_hd__buf_2 _14198_ (.A(_08189_),
    .X(_08207_));
 sky130_fd_sc_hd__nor2_4 _14199_ (.A(\CPU_Xreg_value_a4[15][25] ),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__a211o_4 _14200_ (.A1(_08098_),
    .A2(_08202_),
    .B1(_08198_),
    .C1(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__inv_2 _14201_ (.A(_08209_),
    .Y(_00551_));
 sky130_fd_sc_hd__nor2_4 _14202_ (.A(\CPU_Xreg_value_a4[15][24] ),
    .B(_08207_),
    .Y(_08210_));
 sky130_fd_sc_hd__a211o_4 _14203_ (.A1(_08102_),
    .A2(_08202_),
    .B1(_08198_),
    .C1(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__inv_2 _14204_ (.A(_08211_),
    .Y(_00550_));
 sky130_fd_sc_hd__nor2_4 _14205_ (.A(\CPU_Xreg_value_a4[15][23] ),
    .B(_08207_),
    .Y(_08212_));
 sky130_fd_sc_hd__a211o_4 _14206_ (.A1(_08106_),
    .A2(_08202_),
    .B1(_08198_),
    .C1(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__inv_2 _14207_ (.A(_08213_),
    .Y(_00549_));
 sky130_fd_sc_hd__buf_2 _14208_ (.A(_08128_),
    .X(_08214_));
 sky130_fd_sc_hd__nor2_4 _14209_ (.A(\CPU_Xreg_value_a4[15][22] ),
    .B(_08207_),
    .Y(_08215_));
 sky130_fd_sc_hd__a211o_4 _14210_ (.A1(_08110_),
    .A2(_08202_),
    .B1(_08214_),
    .C1(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__inv_2 _14211_ (.A(_08216_),
    .Y(_00548_));
 sky130_fd_sc_hd__buf_2 _14212_ (.A(_08189_),
    .X(_08217_));
 sky130_fd_sc_hd__nor2_4 _14213_ (.A(\CPU_Xreg_value_a4[15][21] ),
    .B(_08207_),
    .Y(_08218_));
 sky130_fd_sc_hd__a211o_4 _14214_ (.A1(_08113_),
    .A2(_08217_),
    .B1(_08214_),
    .C1(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__inv_2 _14215_ (.A(_08219_),
    .Y(_00547_));
 sky130_fd_sc_hd__nor2_4 _14216_ (.A(\CPU_Xreg_value_a4[15][20] ),
    .B(_08207_),
    .Y(_08220_));
 sky130_fd_sc_hd__a211o_4 _14217_ (.A1(_08116_),
    .A2(_08217_),
    .B1(_08214_),
    .C1(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__inv_2 _14218_ (.A(_08221_),
    .Y(_00546_));
 sky130_fd_sc_hd__buf_2 _14219_ (.A(_08188_),
    .X(_08222_));
 sky130_fd_sc_hd__nor2_4 _14220_ (.A(\CPU_Xreg_value_a4[15][19] ),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__a211o_4 _14221_ (.A1(_08119_),
    .A2(_08217_),
    .B1(_08214_),
    .C1(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__inv_2 _14222_ (.A(_08224_),
    .Y(_00545_));
 sky130_fd_sc_hd__nor2_4 _14223_ (.A(\CPU_Xreg_value_a4[15][18] ),
    .B(_08222_),
    .Y(_08225_));
 sky130_fd_sc_hd__a211o_4 _14224_ (.A1(_08123_),
    .A2(_08217_),
    .B1(_08214_),
    .C1(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__inv_2 _14225_ (.A(_08226_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_4 _14226_ (.A(\CPU_Xreg_value_a4[15][17] ),
    .B(_08222_),
    .Y(_08227_));
 sky130_fd_sc_hd__a211o_4 _14227_ (.A1(_08127_),
    .A2(_08217_),
    .B1(_08214_),
    .C1(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__inv_2 _14228_ (.A(_08228_),
    .Y(_00543_));
 sky130_fd_sc_hd__buf_2 _14229_ (.A(_08128_),
    .X(_08229_));
 sky130_fd_sc_hd__nor2_4 _14230_ (.A(\CPU_Xreg_value_a4[15][16] ),
    .B(_08222_),
    .Y(_08230_));
 sky130_fd_sc_hd__a211o_4 _14231_ (.A1(_08132_),
    .A2(_08217_),
    .B1(_08229_),
    .C1(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__inv_2 _14232_ (.A(_08231_),
    .Y(_00542_));
 sky130_fd_sc_hd__buf_2 _14233_ (.A(_08189_),
    .X(_08232_));
 sky130_fd_sc_hd__nor2_4 _14234_ (.A(\CPU_Xreg_value_a4[15][15] ),
    .B(_08222_),
    .Y(_08233_));
 sky130_fd_sc_hd__a211o_4 _14235_ (.A1(_08135_),
    .A2(_08232_),
    .B1(_08229_),
    .C1(_08233_),
    .X(_08234_));
 sky130_fd_sc_hd__inv_2 _14236_ (.A(_08234_),
    .Y(_00541_));
 sky130_fd_sc_hd__nor2_4 _14237_ (.A(\CPU_Xreg_value_a4[15][14] ),
    .B(_08222_),
    .Y(_08235_));
 sky130_fd_sc_hd__a211o_4 _14238_ (.A1(_08138_),
    .A2(_08232_),
    .B1(_08229_),
    .C1(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__inv_2 _14239_ (.A(_08236_),
    .Y(_00540_));
 sky130_fd_sc_hd__buf_2 _14240_ (.A(_08188_),
    .X(_08237_));
 sky130_fd_sc_hd__nor2_4 _14241_ (.A(\CPU_Xreg_value_a4[15][13] ),
    .B(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__a211o_4 _14242_ (.A1(_08141_),
    .A2(_08232_),
    .B1(_08229_),
    .C1(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__inv_2 _14243_ (.A(_08239_),
    .Y(_00539_));
 sky130_fd_sc_hd__nor2_4 _14244_ (.A(\CPU_Xreg_value_a4[15][12] ),
    .B(_08237_),
    .Y(_08240_));
 sky130_fd_sc_hd__a211o_4 _14245_ (.A1(_08145_),
    .A2(_08232_),
    .B1(_08229_),
    .C1(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__inv_2 _14246_ (.A(_08241_),
    .Y(_00538_));
 sky130_fd_sc_hd__nor2_4 _14247_ (.A(\CPU_Xreg_value_a4[15][11] ),
    .B(_08237_),
    .Y(_08242_));
 sky130_fd_sc_hd__a211o_4 _14248_ (.A1(_08149_),
    .A2(_08232_),
    .B1(_08229_),
    .C1(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__inv_2 _14249_ (.A(_08243_),
    .Y(_00537_));
 sky130_fd_sc_hd__buf_2 _14250_ (.A(_07801_),
    .X(_08244_));
 sky130_fd_sc_hd__buf_2 _14251_ (.A(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__nor2_4 _14252_ (.A(\CPU_Xreg_value_a4[15][10] ),
    .B(_08237_),
    .Y(_08246_));
 sky130_fd_sc_hd__a211o_4 _14253_ (.A1(_08153_),
    .A2(_08232_),
    .B1(_08245_),
    .C1(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__inv_2 _14254_ (.A(_08247_),
    .Y(_00536_));
 sky130_fd_sc_hd__buf_2 _14255_ (.A(_08189_),
    .X(_08248_));
 sky130_fd_sc_hd__nor2_4 _14256_ (.A(\CPU_Xreg_value_a4[15][9] ),
    .B(_08237_),
    .Y(_08249_));
 sky130_fd_sc_hd__a211o_4 _14257_ (.A1(_08156_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__inv_2 _14258_ (.A(_08250_),
    .Y(_00535_));
 sky130_fd_sc_hd__nor2_4 _14259_ (.A(\CPU_Xreg_value_a4[15][8] ),
    .B(_08237_),
    .Y(_08251_));
 sky130_fd_sc_hd__a211o_4 _14260_ (.A1(_08159_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__inv_2 _14261_ (.A(_08252_),
    .Y(_00534_));
 sky130_fd_sc_hd__nor2_4 _14262_ (.A(\CPU_Xreg_value_a4[15][7] ),
    .B(_08201_),
    .Y(_08253_));
 sky130_fd_sc_hd__a211o_4 _14263_ (.A1(_08162_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__inv_2 _14264_ (.A(_08254_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_4 _14265_ (.A(\CPU_Xreg_value_a4[15][6] ),
    .B(_08201_),
    .Y(_08255_));
 sky130_fd_sc_hd__a211o_4 _14266_ (.A1(_08165_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__inv_2 _14267_ (.A(_08256_),
    .Y(_00532_));
 sky130_fd_sc_hd__nor2_4 _14268_ (.A(\CPU_Xreg_value_a4[15][5] ),
    .B(_08201_),
    .Y(_08257_));
 sky130_fd_sc_hd__a211o_4 _14269_ (.A1(_08168_),
    .A2(_08248_),
    .B1(_08245_),
    .C1(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__inv_2 _14270_ (.A(_08258_),
    .Y(_00531_));
 sky130_fd_sc_hd__buf_2 _14271_ (.A(_08244_),
    .X(_08259_));
 sky130_fd_sc_hd__nor2_4 _14272_ (.A(\CPU_Xreg_value_a4[15][4] ),
    .B(_08201_),
    .Y(_08260_));
 sky130_fd_sc_hd__a211o_4 _14273_ (.A1(_06843_),
    .A2(_08248_),
    .B1(_08259_),
    .C1(_08260_),
    .X(_08261_));
 sky130_fd_sc_hd__inv_2 _14274_ (.A(_08261_),
    .Y(_00530_));
 sky130_fd_sc_hd__buf_2 _14275_ (.A(_08201_),
    .X(_08262_));
 sky130_fd_sc_hd__buf_2 _14276_ (.A(_08065_),
    .X(_08263_));
 sky130_fd_sc_hd__inv_2 _14277_ (.A(\CPU_Xreg_value_a4[15][3] ),
    .Y(_08264_));
 sky130_fd_sc_hd__nor2_4 _14278_ (.A(_08264_),
    .B(_08262_),
    .Y(_08265_));
 sky130_fd_sc_hd__a211o_4 _14279_ (.A1(_08174_),
    .A2(_08262_),
    .B1(_08263_),
    .C1(_08265_),
    .X(_00529_));
 sky130_fd_sc_hd__inv_2 _14280_ (.A(\CPU_Xreg_value_a4[15][2] ),
    .Y(_08266_));
 sky130_fd_sc_hd__nor2_4 _14281_ (.A(_08266_),
    .B(_08262_),
    .Y(_08267_));
 sky130_fd_sc_hd__a211o_4 _14282_ (.A1(_08178_),
    .A2(_08262_),
    .B1(_08263_),
    .C1(_08267_),
    .X(_00528_));
 sky130_fd_sc_hd__inv_2 _14283_ (.A(\CPU_Xreg_value_a4[15][1] ),
    .Y(_08268_));
 sky130_fd_sc_hd__nor2_4 _14284_ (.A(_08268_),
    .B(_08190_),
    .Y(_08269_));
 sky130_fd_sc_hd__a211o_4 _14285_ (.A1(_08181_),
    .A2(_08262_),
    .B1(_08263_),
    .C1(_08269_),
    .X(_00527_));
 sky130_fd_sc_hd__buf_2 _14286_ (.A(_06981_),
    .X(_08270_));
 sky130_fd_sc_hd__inv_2 _14287_ (.A(\CPU_Xreg_value_a4[15][0] ),
    .Y(_08271_));
 sky130_fd_sc_hd__nor2_4 _14288_ (.A(_08271_),
    .B(_08190_),
    .Y(_08272_));
 sky130_fd_sc_hd__a211o_4 _14289_ (.A1(_08270_),
    .A2(_08262_),
    .B1(_08263_),
    .C1(_08272_),
    .X(_00526_));
 sky130_fd_sc_hd__or2_4 _14290_ (.A(_06157_),
    .B(_06163_),
    .X(_08273_));
 sky130_fd_sc_hd__inv_2 _14291_ (.A(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__buf_2 _14292_ (.A(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__buf_2 _14293_ (.A(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__buf_2 _14294_ (.A(_08274_),
    .X(_08277_));
 sky130_fd_sc_hd__buf_2 _14295_ (.A(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__nor2_4 _14296_ (.A(\CPU_Xreg_value_a4[16][31] ),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__a211o_4 _14297_ (.A1(_08072_),
    .A2(_08276_),
    .B1(_08259_),
    .C1(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__inv_2 _14298_ (.A(_08280_),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2_4 _14299_ (.A(\CPU_Xreg_value_a4[16][30] ),
    .B(_08278_),
    .Y(_08281_));
 sky130_fd_sc_hd__a211o_4 _14300_ (.A1(_08081_),
    .A2(_08276_),
    .B1(_08259_),
    .C1(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__inv_2 _14301_ (.A(_08282_),
    .Y(_00524_));
 sky130_fd_sc_hd__nor2_4 _14302_ (.A(\CPU_Xreg_value_a4[16][29] ),
    .B(_08278_),
    .Y(_08283_));
 sky130_fd_sc_hd__a211o_4 _14303_ (.A1(_08085_),
    .A2(_08276_),
    .B1(_08259_),
    .C1(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__inv_2 _14304_ (.A(_08284_),
    .Y(_00523_));
 sky130_fd_sc_hd__nor2_4 _14305_ (.A(\CPU_Xreg_value_a4[16][28] ),
    .B(_08278_),
    .Y(_08285_));
 sky130_fd_sc_hd__a211o_4 _14306_ (.A1(_08089_),
    .A2(_08276_),
    .B1(_08259_),
    .C1(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__inv_2 _14307_ (.A(_08286_),
    .Y(_00522_));
 sky130_fd_sc_hd__buf_2 _14308_ (.A(_08277_),
    .X(_08287_));
 sky130_fd_sc_hd__nor2_4 _14309_ (.A(\CPU_Xreg_value_a4[16][27] ),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__a211o_4 _14310_ (.A1(_08092_),
    .A2(_08276_),
    .B1(_08259_),
    .C1(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__inv_2 _14311_ (.A(_08289_),
    .Y(_00521_));
 sky130_fd_sc_hd__buf_2 _14312_ (.A(_08275_),
    .X(_08290_));
 sky130_fd_sc_hd__buf_2 _14313_ (.A(_08244_),
    .X(_08291_));
 sky130_fd_sc_hd__nor2_4 _14314_ (.A(\CPU_Xreg_value_a4[16][26] ),
    .B(_08287_),
    .Y(_08292_));
 sky130_fd_sc_hd__a211o_4 _14315_ (.A1(_08095_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08292_),
    .X(_08293_));
 sky130_fd_sc_hd__inv_2 _14316_ (.A(_08293_),
    .Y(_00520_));
 sky130_fd_sc_hd__nor2_4 _14317_ (.A(\CPU_Xreg_value_a4[16][25] ),
    .B(_08287_),
    .Y(_08294_));
 sky130_fd_sc_hd__a211o_4 _14318_ (.A1(_08098_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__inv_2 _14319_ (.A(_08295_),
    .Y(_00519_));
 sky130_fd_sc_hd__nor2_4 _14320_ (.A(\CPU_Xreg_value_a4[16][24] ),
    .B(_08287_),
    .Y(_08296_));
 sky130_fd_sc_hd__a211o_4 _14321_ (.A1(_08102_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08296_),
    .X(_08297_));
 sky130_fd_sc_hd__inv_2 _14322_ (.A(_08297_),
    .Y(_00518_));
 sky130_fd_sc_hd__nor2_4 _14323_ (.A(\CPU_Xreg_value_a4[16][23] ),
    .B(_08287_),
    .Y(_08298_));
 sky130_fd_sc_hd__a211o_4 _14324_ (.A1(_08106_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__inv_2 _14325_ (.A(_08299_),
    .Y(_00517_));
 sky130_fd_sc_hd__nor2_4 _14326_ (.A(\CPU_Xreg_value_a4[16][22] ),
    .B(_08287_),
    .Y(_08300_));
 sky130_fd_sc_hd__a211o_4 _14327_ (.A1(_08110_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__inv_2 _14328_ (.A(_08301_),
    .Y(_00516_));
 sky130_fd_sc_hd__buf_2 _14329_ (.A(_08277_),
    .X(_08302_));
 sky130_fd_sc_hd__nor2_4 _14330_ (.A(\CPU_Xreg_value_a4[16][21] ),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a211o_4 _14331_ (.A1(_08113_),
    .A2(_08290_),
    .B1(_08291_),
    .C1(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__inv_2 _14332_ (.A(_08304_),
    .Y(_00515_));
 sky130_fd_sc_hd__buf_2 _14333_ (.A(_08275_),
    .X(_08305_));
 sky130_fd_sc_hd__buf_2 _14334_ (.A(_08244_),
    .X(_08306_));
 sky130_fd_sc_hd__nor2_4 _14335_ (.A(\CPU_Xreg_value_a4[16][20] ),
    .B(_08302_),
    .Y(_08307_));
 sky130_fd_sc_hd__a211o_4 _14336_ (.A1(_08116_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__inv_2 _14337_ (.A(_08308_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_4 _14338_ (.A(\CPU_Xreg_value_a4[16][19] ),
    .B(_08302_),
    .Y(_08309_));
 sky130_fd_sc_hd__a211o_4 _14339_ (.A1(_08119_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__inv_2 _14340_ (.A(_08310_),
    .Y(_00513_));
 sky130_fd_sc_hd__nor2_4 _14341_ (.A(\CPU_Xreg_value_a4[16][18] ),
    .B(_08302_),
    .Y(_08311_));
 sky130_fd_sc_hd__a211o_4 _14342_ (.A1(_08123_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__inv_2 _14343_ (.A(_08312_),
    .Y(_00512_));
 sky130_fd_sc_hd__nor2_4 _14344_ (.A(\CPU_Xreg_value_a4[16][17] ),
    .B(_08302_),
    .Y(_08313_));
 sky130_fd_sc_hd__a211o_4 _14345_ (.A1(_08127_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__inv_2 _14346_ (.A(_08314_),
    .Y(_00511_));
 sky130_fd_sc_hd__nor2_4 _14347_ (.A(\CPU_Xreg_value_a4[16][16] ),
    .B(_08302_),
    .Y(_08315_));
 sky130_fd_sc_hd__a211o_4 _14348_ (.A1(_08132_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__inv_2 _14349_ (.A(_08316_),
    .Y(_00510_));
 sky130_fd_sc_hd__buf_2 _14350_ (.A(_08277_),
    .X(_08317_));
 sky130_fd_sc_hd__nor2_4 _14351_ (.A(\CPU_Xreg_value_a4[16][15] ),
    .B(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__a211o_4 _14352_ (.A1(_08135_),
    .A2(_08305_),
    .B1(_08306_),
    .C1(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__inv_2 _14353_ (.A(_08319_),
    .Y(_00509_));
 sky130_fd_sc_hd__buf_2 _14354_ (.A(_08277_),
    .X(_08320_));
 sky130_fd_sc_hd__buf_2 _14355_ (.A(_08244_),
    .X(_08321_));
 sky130_fd_sc_hd__nor2_4 _14356_ (.A(\CPU_Xreg_value_a4[16][14] ),
    .B(_08317_),
    .Y(_08322_));
 sky130_fd_sc_hd__a211o_4 _14357_ (.A1(_08138_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__inv_2 _14358_ (.A(_08323_),
    .Y(_00508_));
 sky130_fd_sc_hd__nor2_4 _14359_ (.A(\CPU_Xreg_value_a4[16][13] ),
    .B(_08317_),
    .Y(_08324_));
 sky130_fd_sc_hd__a211o_4 _14360_ (.A1(_08141_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08324_),
    .X(_08325_));
 sky130_fd_sc_hd__inv_2 _14361_ (.A(_08325_),
    .Y(_00507_));
 sky130_fd_sc_hd__nor2_4 _14362_ (.A(\CPU_Xreg_value_a4[16][12] ),
    .B(_08317_),
    .Y(_08326_));
 sky130_fd_sc_hd__a211o_4 _14363_ (.A1(_08145_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__inv_2 _14364_ (.A(_08327_),
    .Y(_00506_));
 sky130_fd_sc_hd__nor2_4 _14365_ (.A(\CPU_Xreg_value_a4[16][11] ),
    .B(_08317_),
    .Y(_08328_));
 sky130_fd_sc_hd__a211o_4 _14366_ (.A1(_08149_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(_08329_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2_4 _14368_ (.A(\CPU_Xreg_value_a4[16][10] ),
    .B(_08317_),
    .Y(_08330_));
 sky130_fd_sc_hd__a211o_4 _14369_ (.A1(_08153_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__inv_2 _14370_ (.A(_08331_),
    .Y(_00504_));
 sky130_fd_sc_hd__buf_2 _14371_ (.A(_08274_),
    .X(_08332_));
 sky130_fd_sc_hd__nor2_4 _14372_ (.A(\CPU_Xreg_value_a4[16][9] ),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__a211o_4 _14373_ (.A1(_08156_),
    .A2(_08320_),
    .B1(_08321_),
    .C1(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__inv_2 _14374_ (.A(_08334_),
    .Y(_00503_));
 sky130_fd_sc_hd__buf_2 _14375_ (.A(_08277_),
    .X(_08335_));
 sky130_fd_sc_hd__buf_2 _14376_ (.A(_08244_),
    .X(_08336_));
 sky130_fd_sc_hd__nor2_4 _14377_ (.A(\CPU_Xreg_value_a4[16][8] ),
    .B(_08332_),
    .Y(_08337_));
 sky130_fd_sc_hd__a211o_4 _14378_ (.A1(_08159_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__inv_2 _14379_ (.A(_08338_),
    .Y(_00502_));
 sky130_fd_sc_hd__nor2_4 _14380_ (.A(\CPU_Xreg_value_a4[16][7] ),
    .B(_08332_),
    .Y(_08339_));
 sky130_fd_sc_hd__a211o_4 _14381_ (.A1(_08162_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08339_),
    .X(_08340_));
 sky130_fd_sc_hd__inv_2 _14382_ (.A(_08340_),
    .Y(_00501_));
 sky130_fd_sc_hd__nor2_4 _14383_ (.A(\CPU_Xreg_value_a4[16][6] ),
    .B(_08332_),
    .Y(_08341_));
 sky130_fd_sc_hd__a211o_4 _14384_ (.A1(_08165_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__inv_2 _14385_ (.A(_08342_),
    .Y(_00500_));
 sky130_fd_sc_hd__nor2_4 _14386_ (.A(\CPU_Xreg_value_a4[16][5] ),
    .B(_08332_),
    .Y(_08343_));
 sky130_fd_sc_hd__a211o_4 _14387_ (.A1(_08168_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__inv_2 _14388_ (.A(_08344_),
    .Y(_00499_));
 sky130_fd_sc_hd__buf_2 _14389_ (.A(_06842_),
    .X(_08345_));
 sky130_fd_sc_hd__buf_2 _14390_ (.A(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__and2_4 _14391_ (.A(\CPU_Xreg_value_a4[16][4] ),
    .B(_08273_),
    .X(_08347_));
 sky130_fd_sc_hd__a211o_4 _14392_ (.A1(_08346_),
    .A2(_08276_),
    .B1(_08263_),
    .C1(_08347_),
    .X(_00498_));
 sky130_fd_sc_hd__buf_2 _14393_ (.A(_06852_),
    .X(_08348_));
 sky130_fd_sc_hd__nor2_4 _14394_ (.A(\CPU_Xreg_value_a4[16][3] ),
    .B(_08332_),
    .Y(_08349_));
 sky130_fd_sc_hd__a211o_4 _14395_ (.A1(_08348_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__inv_2 _14396_ (.A(_08350_),
    .Y(_00497_));
 sky130_fd_sc_hd__buf_2 _14397_ (.A(_06860_),
    .X(_08351_));
 sky130_fd_sc_hd__nor2_4 _14398_ (.A(\CPU_Xreg_value_a4[16][2] ),
    .B(_08275_),
    .Y(_08352_));
 sky130_fd_sc_hd__a211o_4 _14399_ (.A1(_08351_),
    .A2(_08335_),
    .B1(_08336_),
    .C1(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__inv_2 _14400_ (.A(_08353_),
    .Y(_00496_));
 sky130_fd_sc_hd__buf_2 _14401_ (.A(_06868_),
    .X(_08354_));
 sky130_fd_sc_hd__buf_2 _14402_ (.A(_07801_),
    .X(_08355_));
 sky130_fd_sc_hd__buf_2 _14403_ (.A(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__nor2_4 _14404_ (.A(\CPU_Xreg_value_a4[16][1] ),
    .B(_08275_),
    .Y(_08357_));
 sky130_fd_sc_hd__a211o_4 _14405_ (.A1(_08354_),
    .A2(_08278_),
    .B1(_08356_),
    .C1(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__inv_2 _14406_ (.A(_08358_),
    .Y(_00495_));
 sky130_fd_sc_hd__nor2_4 _14407_ (.A(\CPU_Xreg_value_a4[16][0] ),
    .B(_08275_),
    .Y(_08359_));
 sky130_fd_sc_hd__a211o_4 _14408_ (.A1(_08184_),
    .A2(_08278_),
    .B1(_08356_),
    .C1(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__inv_2 _14409_ (.A(_08360_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_4 _14410_ (.A(_06155_),
    .B(_06162_),
    .Y(_08361_));
 sky130_fd_sc_hd__buf_2 _14411_ (.A(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__buf_2 _14412_ (.A(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__nor2_4 _14413_ (.A(_06153_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__buf_2 _14414_ (.A(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__buf_2 _14415_ (.A(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__buf_2 _14416_ (.A(_08365_),
    .X(_08367_));
 sky130_fd_sc_hd__nor2_4 _14417_ (.A(\CPU_Xreg_value_a4[17][31] ),
    .B(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__a211o_4 _14418_ (.A1(_08072_),
    .A2(_08366_),
    .B1(_08356_),
    .C1(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__inv_2 _14419_ (.A(_08369_),
    .Y(_00493_));
 sky130_fd_sc_hd__nor2_4 _14420_ (.A(\CPU_Xreg_value_a4[17][30] ),
    .B(_08367_),
    .Y(_08370_));
 sky130_fd_sc_hd__a211o_4 _14421_ (.A1(_08081_),
    .A2(_08366_),
    .B1(_08356_),
    .C1(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__inv_2 _14422_ (.A(_08371_),
    .Y(_00492_));
 sky130_fd_sc_hd__buf_2 _14423_ (.A(_08364_),
    .X(_08372_));
 sky130_fd_sc_hd__buf_2 _14424_ (.A(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__buf_2 _14425_ (.A(_08365_),
    .X(_08374_));
 sky130_fd_sc_hd__nor2_4 _14426_ (.A(\CPU_Xreg_value_a4[17][29] ),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__a211o_4 _14427_ (.A1(_08085_),
    .A2(_08373_),
    .B1(_08356_),
    .C1(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__inv_2 _14428_ (.A(_08376_),
    .Y(_00491_));
 sky130_fd_sc_hd__nor2_4 _14429_ (.A(\CPU_Xreg_value_a4[17][28] ),
    .B(_08374_),
    .Y(_08377_));
 sky130_fd_sc_hd__a211o_4 _14430_ (.A1(_08089_),
    .A2(_08373_),
    .B1(_08356_),
    .C1(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__inv_2 _14431_ (.A(_08378_),
    .Y(_00490_));
 sky130_fd_sc_hd__buf_2 _14432_ (.A(_08355_),
    .X(_08379_));
 sky130_fd_sc_hd__nor2_4 _14433_ (.A(\CPU_Xreg_value_a4[17][27] ),
    .B(_08374_),
    .Y(_08380_));
 sky130_fd_sc_hd__a211o_4 _14434_ (.A1(_08092_),
    .A2(_08373_),
    .B1(_08379_),
    .C1(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__inv_2 _14435_ (.A(_08381_),
    .Y(_00489_));
 sky130_fd_sc_hd__nor2_4 _14436_ (.A(\CPU_Xreg_value_a4[17][26] ),
    .B(_08374_),
    .Y(_08382_));
 sky130_fd_sc_hd__a211o_4 _14437_ (.A1(_08095_),
    .A2(_08373_),
    .B1(_08379_),
    .C1(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__inv_2 _14438_ (.A(_08383_),
    .Y(_00488_));
 sky130_fd_sc_hd__nor2_4 _14439_ (.A(\CPU_Xreg_value_a4[17][25] ),
    .B(_08374_),
    .Y(_08384_));
 sky130_fd_sc_hd__a211o_4 _14440_ (.A1(_08098_),
    .A2(_08373_),
    .B1(_08379_),
    .C1(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__inv_2 _14441_ (.A(_08385_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_4 _14442_ (.A(\CPU_Xreg_value_a4[17][24] ),
    .B(_08374_),
    .Y(_08386_));
 sky130_fd_sc_hd__a211o_4 _14443_ (.A1(_08102_),
    .A2(_08373_),
    .B1(_08379_),
    .C1(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__inv_2 _14444_ (.A(_08387_),
    .Y(_00486_));
 sky130_fd_sc_hd__buf_2 _14445_ (.A(_08372_),
    .X(_08388_));
 sky130_fd_sc_hd__buf_2 _14446_ (.A(_08365_),
    .X(_08389_));
 sky130_fd_sc_hd__nor2_4 _14447_ (.A(\CPU_Xreg_value_a4[17][23] ),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__a211o_4 _14448_ (.A1(_08106_),
    .A2(_08388_),
    .B1(_08379_),
    .C1(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__inv_2 _14449_ (.A(_08391_),
    .Y(_00485_));
 sky130_fd_sc_hd__nor2_4 _14450_ (.A(\CPU_Xreg_value_a4[17][22] ),
    .B(_08389_),
    .Y(_08392_));
 sky130_fd_sc_hd__a211o_4 _14451_ (.A1(_08110_),
    .A2(_08388_),
    .B1(_08379_),
    .C1(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__inv_2 _14452_ (.A(_08393_),
    .Y(_00484_));
 sky130_fd_sc_hd__buf_2 _14453_ (.A(_08355_),
    .X(_08394_));
 sky130_fd_sc_hd__nor2_4 _14454_ (.A(\CPU_Xreg_value_a4[17][21] ),
    .B(_08389_),
    .Y(_08395_));
 sky130_fd_sc_hd__a211o_4 _14455_ (.A1(_08113_),
    .A2(_08388_),
    .B1(_08394_),
    .C1(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(_08396_),
    .Y(_00483_));
 sky130_fd_sc_hd__nor2_4 _14457_ (.A(\CPU_Xreg_value_a4[17][20] ),
    .B(_08389_),
    .Y(_08397_));
 sky130_fd_sc_hd__a211o_4 _14458_ (.A1(_08116_),
    .A2(_08388_),
    .B1(_08394_),
    .C1(_08397_),
    .X(_08398_));
 sky130_fd_sc_hd__inv_2 _14459_ (.A(_08398_),
    .Y(_00482_));
 sky130_fd_sc_hd__nor2_4 _14460_ (.A(\CPU_Xreg_value_a4[17][19] ),
    .B(_08389_),
    .Y(_08399_));
 sky130_fd_sc_hd__a211o_4 _14461_ (.A1(_08119_),
    .A2(_08388_),
    .B1(_08394_),
    .C1(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__inv_2 _14462_ (.A(_08400_),
    .Y(_00481_));
 sky130_fd_sc_hd__nor2_4 _14463_ (.A(\CPU_Xreg_value_a4[17][18] ),
    .B(_08389_),
    .Y(_08401_));
 sky130_fd_sc_hd__a211o_4 _14464_ (.A1(_08123_),
    .A2(_08388_),
    .B1(_08394_),
    .C1(_08401_),
    .X(_08402_));
 sky130_fd_sc_hd__inv_2 _14465_ (.A(_08402_),
    .Y(_00480_));
 sky130_fd_sc_hd__buf_2 _14466_ (.A(_08365_),
    .X(_08403_));
 sky130_fd_sc_hd__buf_2 _14467_ (.A(_08364_),
    .X(_08404_));
 sky130_fd_sc_hd__nor2_4 _14468_ (.A(\CPU_Xreg_value_a4[17][17] ),
    .B(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__a211o_4 _14469_ (.A1(_08127_),
    .A2(_08403_),
    .B1(_08394_),
    .C1(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__inv_2 _14470_ (.A(_08406_),
    .Y(_00479_));
 sky130_fd_sc_hd__nor2_4 _14471_ (.A(\CPU_Xreg_value_a4[17][16] ),
    .B(_08404_),
    .Y(_08407_));
 sky130_fd_sc_hd__a211o_4 _14472_ (.A1(_08132_),
    .A2(_08403_),
    .B1(_08394_),
    .C1(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__inv_2 _14473_ (.A(_08408_),
    .Y(_00478_));
 sky130_fd_sc_hd__buf_2 _14474_ (.A(_08355_),
    .X(_08409_));
 sky130_fd_sc_hd__nor2_4 _14475_ (.A(\CPU_Xreg_value_a4[17][15] ),
    .B(_08404_),
    .Y(_08410_));
 sky130_fd_sc_hd__a211o_4 _14476_ (.A1(_08135_),
    .A2(_08403_),
    .B1(_08409_),
    .C1(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__inv_2 _14477_ (.A(_08411_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_4 _14478_ (.A(\CPU_Xreg_value_a4[17][14] ),
    .B(_08404_),
    .Y(_08412_));
 sky130_fd_sc_hd__a211o_4 _14479_ (.A1(_08138_),
    .A2(_08403_),
    .B1(_08409_),
    .C1(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__inv_2 _14480_ (.A(_08413_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_4 _14481_ (.A(\CPU_Xreg_value_a4[17][13] ),
    .B(_08404_),
    .Y(_08414_));
 sky130_fd_sc_hd__a211o_4 _14482_ (.A1(_08141_),
    .A2(_08403_),
    .B1(_08409_),
    .C1(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__inv_2 _14483_ (.A(_08415_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_4 _14484_ (.A(\CPU_Xreg_value_a4[17][12] ),
    .B(_08404_),
    .Y(_08416_));
 sky130_fd_sc_hd__a211o_4 _14485_ (.A1(_08145_),
    .A2(_08403_),
    .B1(_08409_),
    .C1(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__inv_2 _14486_ (.A(_08417_),
    .Y(_00474_));
 sky130_fd_sc_hd__buf_2 _14487_ (.A(_08365_),
    .X(_08418_));
 sky130_fd_sc_hd__buf_2 _14488_ (.A(_08364_),
    .X(_08419_));
 sky130_fd_sc_hd__nor2_4 _14489_ (.A(\CPU_Xreg_value_a4[17][11] ),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__a211o_4 _14490_ (.A1(_08149_),
    .A2(_08418_),
    .B1(_08409_),
    .C1(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__inv_2 _14491_ (.A(_08421_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_4 _14492_ (.A(\CPU_Xreg_value_a4[17][10] ),
    .B(_08419_),
    .Y(_08422_));
 sky130_fd_sc_hd__a211o_4 _14493_ (.A1(_08153_),
    .A2(_08418_),
    .B1(_08409_),
    .C1(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__inv_2 _14494_ (.A(_08423_),
    .Y(_00472_));
 sky130_fd_sc_hd__buf_2 _14495_ (.A(_08355_),
    .X(_08424_));
 sky130_fd_sc_hd__nor2_4 _14496_ (.A(\CPU_Xreg_value_a4[17][9] ),
    .B(_08419_),
    .Y(_08425_));
 sky130_fd_sc_hd__a211o_4 _14497_ (.A1(_08156_),
    .A2(_08418_),
    .B1(_08424_),
    .C1(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__inv_2 _14498_ (.A(_08426_),
    .Y(_00471_));
 sky130_fd_sc_hd__nor2_4 _14499_ (.A(\CPU_Xreg_value_a4[17][8] ),
    .B(_08419_),
    .Y(_08427_));
 sky130_fd_sc_hd__a211o_4 _14500_ (.A1(_08159_),
    .A2(_08418_),
    .B1(_08424_),
    .C1(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__inv_2 _14501_ (.A(_08428_),
    .Y(_00470_));
 sky130_fd_sc_hd__nor2_4 _14502_ (.A(\CPU_Xreg_value_a4[17][7] ),
    .B(_08419_),
    .Y(_08429_));
 sky130_fd_sc_hd__a211o_4 _14503_ (.A1(_08162_),
    .A2(_08418_),
    .B1(_08424_),
    .C1(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__inv_2 _14504_ (.A(_08430_),
    .Y(_00469_));
 sky130_fd_sc_hd__nor2_4 _14505_ (.A(\CPU_Xreg_value_a4[17][6] ),
    .B(_08419_),
    .Y(_08431_));
 sky130_fd_sc_hd__a211o_4 _14506_ (.A1(_08165_),
    .A2(_08418_),
    .B1(_08424_),
    .C1(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__inv_2 _14507_ (.A(_08432_),
    .Y(_00468_));
 sky130_fd_sc_hd__nor2_4 _14508_ (.A(\CPU_Xreg_value_a4[17][5] ),
    .B(_08372_),
    .Y(_08433_));
 sky130_fd_sc_hd__a211o_4 _14509_ (.A1(_08168_),
    .A2(_08367_),
    .B1(_08424_),
    .C1(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__inv_2 _14510_ (.A(_08434_),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _14511_ (.A(\CPU_Xreg_value_a4[17][4] ),
    .Y(_08435_));
 sky130_fd_sc_hd__nor2_4 _14512_ (.A(_08435_),
    .B(_08366_),
    .Y(_08436_));
 sky130_fd_sc_hd__a211o_4 _14513_ (.A1(_08346_),
    .A2(_08366_),
    .B1(_08263_),
    .C1(_08436_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_4 _14514_ (.A(\CPU_Xreg_value_a4[17][3] ),
    .B(_08372_),
    .Y(_08437_));
 sky130_fd_sc_hd__a211o_4 _14515_ (.A1(_08348_),
    .A2(_08367_),
    .B1(_08424_),
    .C1(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__inv_2 _14516_ (.A(_08438_),
    .Y(_00465_));
 sky130_fd_sc_hd__buf_2 _14517_ (.A(_08355_),
    .X(_08439_));
 sky130_fd_sc_hd__nor2_4 _14518_ (.A(\CPU_Xreg_value_a4[17][2] ),
    .B(_08372_),
    .Y(_08440_));
 sky130_fd_sc_hd__a211o_4 _14519_ (.A1(_08351_),
    .A2(_08367_),
    .B1(_08439_),
    .C1(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__inv_2 _14520_ (.A(_08441_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_4 _14521_ (.A(\CPU_Xreg_value_a4[17][1] ),
    .B(_08372_),
    .Y(_08442_));
 sky130_fd_sc_hd__a211o_4 _14522_ (.A1(_08354_),
    .A2(_08367_),
    .B1(_08439_),
    .C1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__inv_2 _14523_ (.A(_08443_),
    .Y(_00463_));
 sky130_fd_sc_hd__buf_2 _14524_ (.A(_08065_),
    .X(_08444_));
 sky130_fd_sc_hd__inv_2 _14525_ (.A(\CPU_Xreg_value_a4[17][0] ),
    .Y(_08445_));
 sky130_fd_sc_hd__nor2_4 _14526_ (.A(_08445_),
    .B(_08366_),
    .Y(_08446_));
 sky130_fd_sc_hd__a211o_4 _14527_ (.A1(_08270_),
    .A2(_08366_),
    .B1(_08444_),
    .C1(_08446_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_4 _14528_ (.A(_06987_),
    .B(_08363_),
    .Y(_08447_));
 sky130_fd_sc_hd__buf_2 _14529_ (.A(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__buf_2 _14530_ (.A(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__buf_2 _14531_ (.A(_08448_),
    .X(_08450_));
 sky130_fd_sc_hd__nor2_4 _14532_ (.A(\CPU_Xreg_value_a4[18][31] ),
    .B(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__a211o_4 _14533_ (.A1(_08072_),
    .A2(_08449_),
    .B1(_08439_),
    .C1(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__inv_2 _14534_ (.A(_08452_),
    .Y(_00461_));
 sky130_fd_sc_hd__nor2_4 _14535_ (.A(\CPU_Xreg_value_a4[18][30] ),
    .B(_08450_),
    .Y(_08453_));
 sky130_fd_sc_hd__a211o_4 _14536_ (.A1(_08081_),
    .A2(_08449_),
    .B1(_08439_),
    .C1(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__inv_2 _14537_ (.A(_08454_),
    .Y(_00460_));
 sky130_fd_sc_hd__buf_2 _14538_ (.A(_08447_),
    .X(_08455_));
 sky130_fd_sc_hd__buf_2 _14539_ (.A(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__buf_2 _14540_ (.A(_08448_),
    .X(_08457_));
 sky130_fd_sc_hd__nor2_4 _14541_ (.A(\CPU_Xreg_value_a4[18][29] ),
    .B(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__a211o_4 _14542_ (.A1(_08085_),
    .A2(_08456_),
    .B1(_08439_),
    .C1(_08458_),
    .X(_08459_));
 sky130_fd_sc_hd__inv_2 _14543_ (.A(_08459_),
    .Y(_00459_));
 sky130_fd_sc_hd__nor2_4 _14544_ (.A(\CPU_Xreg_value_a4[18][28] ),
    .B(_08457_),
    .Y(_08460_));
 sky130_fd_sc_hd__a211o_4 _14545_ (.A1(_08089_),
    .A2(_08456_),
    .B1(_08439_),
    .C1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__inv_2 _14546_ (.A(_08461_),
    .Y(_00458_));
 sky130_fd_sc_hd__buf_2 _14547_ (.A(CPU_reset_a3),
    .X(_08462_));
 sky130_fd_sc_hd__buf_2 _14548_ (.A(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__buf_2 _14549_ (.A(_08463_),
    .X(_08464_));
 sky130_fd_sc_hd__nor2_4 _14550_ (.A(\CPU_Xreg_value_a4[18][27] ),
    .B(_08457_),
    .Y(_08465_));
 sky130_fd_sc_hd__a211o_4 _14551_ (.A1(_08092_),
    .A2(_08456_),
    .B1(_08464_),
    .C1(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__inv_2 _14552_ (.A(_08466_),
    .Y(_00457_));
 sky130_fd_sc_hd__nor2_4 _14553_ (.A(\CPU_Xreg_value_a4[18][26] ),
    .B(_08457_),
    .Y(_08467_));
 sky130_fd_sc_hd__a211o_4 _14554_ (.A1(_08095_),
    .A2(_08456_),
    .B1(_08464_),
    .C1(_08467_),
    .X(_08468_));
 sky130_fd_sc_hd__inv_2 _14555_ (.A(_08468_),
    .Y(_00456_));
 sky130_fd_sc_hd__nor2_4 _14556_ (.A(\CPU_Xreg_value_a4[18][25] ),
    .B(_08457_),
    .Y(_08469_));
 sky130_fd_sc_hd__a211o_4 _14557_ (.A1(_08098_),
    .A2(_08456_),
    .B1(_08464_),
    .C1(_08469_),
    .X(_08470_));
 sky130_fd_sc_hd__inv_2 _14558_ (.A(_08470_),
    .Y(_00455_));
 sky130_fd_sc_hd__nor2_4 _14559_ (.A(\CPU_Xreg_value_a4[18][24] ),
    .B(_08457_),
    .Y(_08471_));
 sky130_fd_sc_hd__a211o_4 _14560_ (.A1(_08102_),
    .A2(_08456_),
    .B1(_08464_),
    .C1(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__inv_2 _14561_ (.A(_08472_),
    .Y(_00454_));
 sky130_fd_sc_hd__buf_2 _14562_ (.A(_08455_),
    .X(_08473_));
 sky130_fd_sc_hd__buf_2 _14563_ (.A(_08448_),
    .X(_08474_));
 sky130_fd_sc_hd__nor2_4 _14564_ (.A(\CPU_Xreg_value_a4[18][23] ),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__a211o_4 _14565_ (.A1(_08106_),
    .A2(_08473_),
    .B1(_08464_),
    .C1(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__inv_2 _14566_ (.A(_08476_),
    .Y(_00453_));
 sky130_fd_sc_hd__nor2_4 _14567_ (.A(\CPU_Xreg_value_a4[18][22] ),
    .B(_08474_),
    .Y(_08477_));
 sky130_fd_sc_hd__a211o_4 _14568_ (.A1(_08110_),
    .A2(_08473_),
    .B1(_08464_),
    .C1(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__inv_2 _14569_ (.A(_08478_),
    .Y(_00452_));
 sky130_fd_sc_hd__buf_2 _14570_ (.A(_08463_),
    .X(_08479_));
 sky130_fd_sc_hd__nor2_4 _14571_ (.A(\CPU_Xreg_value_a4[18][21] ),
    .B(_08474_),
    .Y(_08480_));
 sky130_fd_sc_hd__a211o_4 _14572_ (.A1(_08113_),
    .A2(_08473_),
    .B1(_08479_),
    .C1(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__inv_2 _14573_ (.A(_08481_),
    .Y(_00451_));
 sky130_fd_sc_hd__nor2_4 _14574_ (.A(\CPU_Xreg_value_a4[18][20] ),
    .B(_08474_),
    .Y(_08482_));
 sky130_fd_sc_hd__a211o_4 _14575_ (.A1(_08116_),
    .A2(_08473_),
    .B1(_08479_),
    .C1(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__inv_2 _14576_ (.A(_08483_),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_4 _14577_ (.A(\CPU_Xreg_value_a4[18][19] ),
    .B(_08474_),
    .Y(_08484_));
 sky130_fd_sc_hd__a211o_4 _14578_ (.A1(_08119_),
    .A2(_08473_),
    .B1(_08479_),
    .C1(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__inv_2 _14579_ (.A(_08485_),
    .Y(_00449_));
 sky130_fd_sc_hd__nor2_4 _14580_ (.A(\CPU_Xreg_value_a4[18][18] ),
    .B(_08474_),
    .Y(_08486_));
 sky130_fd_sc_hd__a211o_4 _14581_ (.A1(_08123_),
    .A2(_08473_),
    .B1(_08479_),
    .C1(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__inv_2 _14582_ (.A(_08487_),
    .Y(_00448_));
 sky130_fd_sc_hd__buf_2 _14583_ (.A(_08448_),
    .X(_08488_));
 sky130_fd_sc_hd__buf_2 _14584_ (.A(_08447_),
    .X(_08489_));
 sky130_fd_sc_hd__nor2_4 _14585_ (.A(\CPU_Xreg_value_a4[18][17] ),
    .B(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__a211o_4 _14586_ (.A1(_08127_),
    .A2(_08488_),
    .B1(_08479_),
    .C1(_08490_),
    .X(_08491_));
 sky130_fd_sc_hd__inv_2 _14587_ (.A(_08491_),
    .Y(_00447_));
 sky130_fd_sc_hd__nor2_4 _14588_ (.A(\CPU_Xreg_value_a4[18][16] ),
    .B(_08489_),
    .Y(_08492_));
 sky130_fd_sc_hd__a211o_4 _14589_ (.A1(_08132_),
    .A2(_08488_),
    .B1(_08479_),
    .C1(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__inv_2 _14590_ (.A(_08493_),
    .Y(_00446_));
 sky130_fd_sc_hd__buf_2 _14591_ (.A(_08463_),
    .X(_08494_));
 sky130_fd_sc_hd__nor2_4 _14592_ (.A(\CPU_Xreg_value_a4[18][15] ),
    .B(_08489_),
    .Y(_08495_));
 sky130_fd_sc_hd__a211o_4 _14593_ (.A1(_08135_),
    .A2(_08488_),
    .B1(_08494_),
    .C1(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__inv_2 _14594_ (.A(_08496_),
    .Y(_00445_));
 sky130_fd_sc_hd__nor2_4 _14595_ (.A(\CPU_Xreg_value_a4[18][14] ),
    .B(_08489_),
    .Y(_08497_));
 sky130_fd_sc_hd__a211o_4 _14596_ (.A1(_08138_),
    .A2(_08488_),
    .B1(_08494_),
    .C1(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__inv_2 _14597_ (.A(_08498_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_4 _14598_ (.A(\CPU_Xreg_value_a4[18][13] ),
    .B(_08489_),
    .Y(_08499_));
 sky130_fd_sc_hd__a211o_4 _14599_ (.A1(_08141_),
    .A2(_08488_),
    .B1(_08494_),
    .C1(_08499_),
    .X(_08500_));
 sky130_fd_sc_hd__inv_2 _14600_ (.A(_08500_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor2_4 _14601_ (.A(\CPU_Xreg_value_a4[18][12] ),
    .B(_08489_),
    .Y(_08501_));
 sky130_fd_sc_hd__a211o_4 _14602_ (.A1(_08145_),
    .A2(_08488_),
    .B1(_08494_),
    .C1(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__inv_2 _14603_ (.A(_08502_),
    .Y(_00442_));
 sky130_fd_sc_hd__buf_2 _14604_ (.A(_08448_),
    .X(_08503_));
 sky130_fd_sc_hd__buf_2 _14605_ (.A(_08447_),
    .X(_08504_));
 sky130_fd_sc_hd__nor2_4 _14606_ (.A(\CPU_Xreg_value_a4[18][11] ),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__a211o_4 _14607_ (.A1(_08149_),
    .A2(_08503_),
    .B1(_08494_),
    .C1(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__inv_2 _14608_ (.A(_08506_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2_4 _14609_ (.A(\CPU_Xreg_value_a4[18][10] ),
    .B(_08504_),
    .Y(_08507_));
 sky130_fd_sc_hd__a211o_4 _14610_ (.A1(_08153_),
    .A2(_08503_),
    .B1(_08494_),
    .C1(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__inv_2 _14611_ (.A(_08508_),
    .Y(_00440_));
 sky130_fd_sc_hd__buf_2 _14612_ (.A(_08463_),
    .X(_08509_));
 sky130_fd_sc_hd__nor2_4 _14613_ (.A(\CPU_Xreg_value_a4[18][9] ),
    .B(_08504_),
    .Y(_08510_));
 sky130_fd_sc_hd__a211o_4 _14614_ (.A1(_08156_),
    .A2(_08503_),
    .B1(_08509_),
    .C1(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__inv_2 _14615_ (.A(_08511_),
    .Y(_00439_));
 sky130_fd_sc_hd__nor2_4 _14616_ (.A(\CPU_Xreg_value_a4[18][8] ),
    .B(_08504_),
    .Y(_08512_));
 sky130_fd_sc_hd__a211o_4 _14617_ (.A1(_08159_),
    .A2(_08503_),
    .B1(_08509_),
    .C1(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__inv_2 _14618_ (.A(_08513_),
    .Y(_00438_));
 sky130_fd_sc_hd__nor2_4 _14619_ (.A(\CPU_Xreg_value_a4[18][7] ),
    .B(_08504_),
    .Y(_08514_));
 sky130_fd_sc_hd__a211o_4 _14620_ (.A1(_08162_),
    .A2(_08503_),
    .B1(_08509_),
    .C1(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__inv_2 _14621_ (.A(_08515_),
    .Y(_00437_));
 sky130_fd_sc_hd__nor2_4 _14622_ (.A(\CPU_Xreg_value_a4[18][6] ),
    .B(_08504_),
    .Y(_08516_));
 sky130_fd_sc_hd__a211o_4 _14623_ (.A1(_08165_),
    .A2(_08503_),
    .B1(_08509_),
    .C1(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__inv_2 _14624_ (.A(_08517_),
    .Y(_00436_));
 sky130_fd_sc_hd__nor2_4 _14625_ (.A(\CPU_Xreg_value_a4[18][5] ),
    .B(_08455_),
    .Y(_08518_));
 sky130_fd_sc_hd__a211o_4 _14626_ (.A1(_08168_),
    .A2(_08450_),
    .B1(_08509_),
    .C1(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__inv_2 _14627_ (.A(_08519_),
    .Y(_00435_));
 sky130_fd_sc_hd__inv_2 _14628_ (.A(\CPU_Xreg_value_a4[18][4] ),
    .Y(_08520_));
 sky130_fd_sc_hd__nor2_4 _14629_ (.A(_08520_),
    .B(_08449_),
    .Y(_08521_));
 sky130_fd_sc_hd__a211o_4 _14630_ (.A1(_08346_),
    .A2(_08449_),
    .B1(_08444_),
    .C1(_08521_),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_4 _14631_ (.A(\CPU_Xreg_value_a4[18][3] ),
    .B(_08455_),
    .Y(_08522_));
 sky130_fd_sc_hd__a211o_4 _14632_ (.A1(_08348_),
    .A2(_08450_),
    .B1(_08509_),
    .C1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__inv_2 _14633_ (.A(_08523_),
    .Y(_00433_));
 sky130_fd_sc_hd__buf_2 _14634_ (.A(_08463_),
    .X(_08524_));
 sky130_fd_sc_hd__nor2_4 _14635_ (.A(\CPU_Xreg_value_a4[18][2] ),
    .B(_08455_),
    .Y(_08525_));
 sky130_fd_sc_hd__a211o_4 _14636_ (.A1(_08351_),
    .A2(_08450_),
    .B1(_08524_),
    .C1(_08525_),
    .X(_08526_));
 sky130_fd_sc_hd__inv_2 _14637_ (.A(_08526_),
    .Y(_00432_));
 sky130_fd_sc_hd__inv_2 _14638_ (.A(\CPU_Xreg_value_a4[18][1] ),
    .Y(_08527_));
 sky130_fd_sc_hd__nor2_4 _14639_ (.A(_08527_),
    .B(_08449_),
    .Y(_08528_));
 sky130_fd_sc_hd__a211o_4 _14640_ (.A1(_08181_),
    .A2(_08449_),
    .B1(_08444_),
    .C1(_08528_),
    .X(_00431_));
 sky130_fd_sc_hd__nor2_4 _14641_ (.A(\CPU_Xreg_value_a4[18][0] ),
    .B(_08455_),
    .Y(_08529_));
 sky130_fd_sc_hd__a211o_4 _14642_ (.A1(_08184_),
    .A2(_08450_),
    .B1(_08524_),
    .C1(_08529_),
    .X(_08530_));
 sky130_fd_sc_hd__inv_2 _14643_ (.A(_08530_),
    .Y(_00430_));
 sky130_fd_sc_hd__nor2_4 _14644_ (.A(_07105_),
    .B(_08363_),
    .Y(_08531_));
 sky130_fd_sc_hd__buf_2 _14645_ (.A(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__buf_2 _14646_ (.A(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__buf_2 _14647_ (.A(_08531_),
    .X(_08534_));
 sky130_fd_sc_hd__buf_2 _14648_ (.A(_08534_),
    .X(_08535_));
 sky130_fd_sc_hd__nor2_4 _14649_ (.A(\CPU_Xreg_value_a4[19][31] ),
    .B(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__a211o_4 _14650_ (.A1(_08072_),
    .A2(_08533_),
    .B1(_08524_),
    .C1(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__inv_2 _14651_ (.A(_08537_),
    .Y(_00429_));
 sky130_fd_sc_hd__buf_2 _14652_ (.A(_08534_),
    .X(_08538_));
 sky130_fd_sc_hd__nor2_4 _14653_ (.A(\CPU_Xreg_value_a4[19][30] ),
    .B(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__a211o_4 _14654_ (.A1(_08081_),
    .A2(_08533_),
    .B1(_08524_),
    .C1(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__inv_2 _14655_ (.A(_08540_),
    .Y(_00428_));
 sky130_fd_sc_hd__nor2_4 _14656_ (.A(\CPU_Xreg_value_a4[19][29] ),
    .B(_08538_),
    .Y(_08541_));
 sky130_fd_sc_hd__a211o_4 _14657_ (.A1(_08085_),
    .A2(_08533_),
    .B1(_08524_),
    .C1(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__inv_2 _14658_ (.A(_08542_),
    .Y(_00427_));
 sky130_fd_sc_hd__nor2_4 _14659_ (.A(\CPU_Xreg_value_a4[19][28] ),
    .B(_08538_),
    .Y(_08543_));
 sky130_fd_sc_hd__a211o_4 _14660_ (.A1(_08089_),
    .A2(_08533_),
    .B1(_08524_),
    .C1(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__inv_2 _14661_ (.A(_08544_),
    .Y(_00426_));
 sky130_fd_sc_hd__buf_2 _14662_ (.A(_08463_),
    .X(_08545_));
 sky130_fd_sc_hd__nor2_4 _14663_ (.A(\CPU_Xreg_value_a4[19][27] ),
    .B(_08538_),
    .Y(_08546_));
 sky130_fd_sc_hd__a211o_4 _14664_ (.A1(_08092_),
    .A2(_08533_),
    .B1(_08545_),
    .C1(_08546_),
    .X(_08547_));
 sky130_fd_sc_hd__inv_2 _14665_ (.A(_08547_),
    .Y(_00425_));
 sky130_fd_sc_hd__nor2_4 _14666_ (.A(\CPU_Xreg_value_a4[19][26] ),
    .B(_08538_),
    .Y(_08548_));
 sky130_fd_sc_hd__a211o_4 _14667_ (.A1(_08095_),
    .A2(_08533_),
    .B1(_08545_),
    .C1(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__inv_2 _14668_ (.A(_08549_),
    .Y(_00424_));
 sky130_fd_sc_hd__buf_2 _14669_ (.A(_08534_),
    .X(_08550_));
 sky130_fd_sc_hd__nor2_4 _14670_ (.A(\CPU_Xreg_value_a4[19][25] ),
    .B(_08538_),
    .Y(_08551_));
 sky130_fd_sc_hd__a211o_4 _14671_ (.A1(_08098_),
    .A2(_08550_),
    .B1(_08545_),
    .C1(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__inv_2 _14672_ (.A(_08552_),
    .Y(_00423_));
 sky130_fd_sc_hd__buf_2 _14673_ (.A(_08534_),
    .X(_08553_));
 sky130_fd_sc_hd__nor2_4 _14674_ (.A(\CPU_Xreg_value_a4[19][24] ),
    .B(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__a211o_4 _14675_ (.A1(_08102_),
    .A2(_08550_),
    .B1(_08545_),
    .C1(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__inv_2 _14676_ (.A(_08555_),
    .Y(_00422_));
 sky130_fd_sc_hd__nor2_4 _14677_ (.A(\CPU_Xreg_value_a4[19][23] ),
    .B(_08553_),
    .Y(_08556_));
 sky130_fd_sc_hd__a211o_4 _14678_ (.A1(_08106_),
    .A2(_08550_),
    .B1(_08545_),
    .C1(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__inv_2 _14679_ (.A(_08557_),
    .Y(_00421_));
 sky130_fd_sc_hd__nor2_4 _14680_ (.A(\CPU_Xreg_value_a4[19][22] ),
    .B(_08553_),
    .Y(_08558_));
 sky130_fd_sc_hd__a211o_4 _14681_ (.A1(_08110_),
    .A2(_08550_),
    .B1(_08545_),
    .C1(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__inv_2 _14682_ (.A(_08559_),
    .Y(_00420_));
 sky130_fd_sc_hd__buf_2 _14683_ (.A(_08462_),
    .X(_08560_));
 sky130_fd_sc_hd__buf_2 _14684_ (.A(_08560_),
    .X(_08561_));
 sky130_fd_sc_hd__nor2_4 _14685_ (.A(\CPU_Xreg_value_a4[19][21] ),
    .B(_08553_),
    .Y(_08562_));
 sky130_fd_sc_hd__a211o_4 _14686_ (.A1(_08113_),
    .A2(_08550_),
    .B1(_08561_),
    .C1(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__inv_2 _14687_ (.A(_08563_),
    .Y(_00419_));
 sky130_fd_sc_hd__nor2_4 _14688_ (.A(\CPU_Xreg_value_a4[19][20] ),
    .B(_08553_),
    .Y(_08564_));
 sky130_fd_sc_hd__a211o_4 _14689_ (.A1(_08116_),
    .A2(_08550_),
    .B1(_08561_),
    .C1(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__inv_2 _14690_ (.A(_08565_),
    .Y(_00418_));
 sky130_fd_sc_hd__buf_2 _14691_ (.A(_08534_),
    .X(_08566_));
 sky130_fd_sc_hd__nor2_4 _14692_ (.A(\CPU_Xreg_value_a4[19][19] ),
    .B(_08553_),
    .Y(_08567_));
 sky130_fd_sc_hd__a211o_4 _14693_ (.A1(_08119_),
    .A2(_08566_),
    .B1(_08561_),
    .C1(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__inv_2 _14694_ (.A(_08568_),
    .Y(_00417_));
 sky130_fd_sc_hd__buf_2 _14695_ (.A(_08531_),
    .X(_08569_));
 sky130_fd_sc_hd__nor2_4 _14696_ (.A(\CPU_Xreg_value_a4[19][18] ),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__a211o_4 _14697_ (.A1(_08123_),
    .A2(_08566_),
    .B1(_08561_),
    .C1(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__inv_2 _14698_ (.A(_08571_),
    .Y(_00416_));
 sky130_fd_sc_hd__nor2_4 _14699_ (.A(\CPU_Xreg_value_a4[19][17] ),
    .B(_08569_),
    .Y(_08572_));
 sky130_fd_sc_hd__a211o_4 _14700_ (.A1(_08127_),
    .A2(_08566_),
    .B1(_08561_),
    .C1(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__inv_2 _14701_ (.A(_08573_),
    .Y(_00415_));
 sky130_fd_sc_hd__nor2_4 _14702_ (.A(\CPU_Xreg_value_a4[19][16] ),
    .B(_08569_),
    .Y(_08574_));
 sky130_fd_sc_hd__a211o_4 _14703_ (.A1(_08132_),
    .A2(_08566_),
    .B1(_08561_),
    .C1(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__inv_2 _14704_ (.A(_08575_),
    .Y(_00414_));
 sky130_fd_sc_hd__buf_2 _14705_ (.A(_08560_),
    .X(_08576_));
 sky130_fd_sc_hd__nor2_4 _14706_ (.A(\CPU_Xreg_value_a4[19][15] ),
    .B(_08569_),
    .Y(_08577_));
 sky130_fd_sc_hd__a211o_4 _14707_ (.A1(_08135_),
    .A2(_08566_),
    .B1(_08576_),
    .C1(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__inv_2 _14708_ (.A(_08578_),
    .Y(_00413_));
 sky130_fd_sc_hd__nor2_4 _14709_ (.A(\CPU_Xreg_value_a4[19][14] ),
    .B(_08569_),
    .Y(_08579_));
 sky130_fd_sc_hd__a211o_4 _14710_ (.A1(_08138_),
    .A2(_08566_),
    .B1(_08576_),
    .C1(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__inv_2 _14711_ (.A(_08580_),
    .Y(_00412_));
 sky130_fd_sc_hd__buf_2 _14712_ (.A(_08534_),
    .X(_08581_));
 sky130_fd_sc_hd__nor2_4 _14713_ (.A(\CPU_Xreg_value_a4[19][13] ),
    .B(_08569_),
    .Y(_08582_));
 sky130_fd_sc_hd__a211o_4 _14714_ (.A1(_08141_),
    .A2(_08581_),
    .B1(_08576_),
    .C1(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__inv_2 _14715_ (.A(_08583_),
    .Y(_00411_));
 sky130_fd_sc_hd__buf_2 _14716_ (.A(_08531_),
    .X(_08584_));
 sky130_fd_sc_hd__nor2_4 _14717_ (.A(\CPU_Xreg_value_a4[19][12] ),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__a211o_4 _14718_ (.A1(_08145_),
    .A2(_08581_),
    .B1(_08576_),
    .C1(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__inv_2 _14719_ (.A(_08586_),
    .Y(_00410_));
 sky130_fd_sc_hd__nor2_4 _14720_ (.A(\CPU_Xreg_value_a4[19][11] ),
    .B(_08584_),
    .Y(_08587_));
 sky130_fd_sc_hd__a211o_4 _14721_ (.A1(_08149_),
    .A2(_08581_),
    .B1(_08576_),
    .C1(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__inv_2 _14722_ (.A(_08588_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2_4 _14723_ (.A(\CPU_Xreg_value_a4[19][10] ),
    .B(_08584_),
    .Y(_08589_));
 sky130_fd_sc_hd__a211o_4 _14724_ (.A1(_08153_),
    .A2(_08581_),
    .B1(_08576_),
    .C1(_08589_),
    .X(_08590_));
 sky130_fd_sc_hd__inv_2 _14725_ (.A(_08590_),
    .Y(_00408_));
 sky130_fd_sc_hd__buf_2 _14726_ (.A(_08560_),
    .X(_08591_));
 sky130_fd_sc_hd__nor2_4 _14727_ (.A(\CPU_Xreg_value_a4[19][9] ),
    .B(_08584_),
    .Y(_08592_));
 sky130_fd_sc_hd__a211o_4 _14728_ (.A1(_08156_),
    .A2(_08581_),
    .B1(_08591_),
    .C1(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__inv_2 _14729_ (.A(_08593_),
    .Y(_00407_));
 sky130_fd_sc_hd__nor2_4 _14730_ (.A(\CPU_Xreg_value_a4[19][8] ),
    .B(_08584_),
    .Y(_08594_));
 sky130_fd_sc_hd__a211o_4 _14731_ (.A1(_08159_),
    .A2(_08581_),
    .B1(_08591_),
    .C1(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__inv_2 _14732_ (.A(_08595_),
    .Y(_00406_));
 sky130_fd_sc_hd__nor2_4 _14733_ (.A(\CPU_Xreg_value_a4[19][7] ),
    .B(_08584_),
    .Y(_08596_));
 sky130_fd_sc_hd__a211o_4 _14734_ (.A1(_08162_),
    .A2(_08535_),
    .B1(_08591_),
    .C1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__inv_2 _14735_ (.A(_08597_),
    .Y(_00405_));
 sky130_fd_sc_hd__nor2_4 _14736_ (.A(\CPU_Xreg_value_a4[19][6] ),
    .B(_08532_),
    .Y(_08598_));
 sky130_fd_sc_hd__a211o_4 _14737_ (.A1(_08165_),
    .A2(_08535_),
    .B1(_08591_),
    .C1(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__inv_2 _14738_ (.A(_08599_),
    .Y(_00404_));
 sky130_fd_sc_hd__nor2_4 _14739_ (.A(\CPU_Xreg_value_a4[19][5] ),
    .B(_08532_),
    .Y(_08600_));
 sky130_fd_sc_hd__a211o_4 _14740_ (.A1(_08168_),
    .A2(_08535_),
    .B1(_08591_),
    .C1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__inv_2 _14741_ (.A(_08601_),
    .Y(_00403_));
 sky130_fd_sc_hd__buf_2 _14742_ (.A(_08532_),
    .X(_08602_));
 sky130_fd_sc_hd__inv_2 _14743_ (.A(\CPU_Xreg_value_a4[19][4] ),
    .Y(_08603_));
 sky130_fd_sc_hd__nor2_4 _14744_ (.A(_08603_),
    .B(_08602_),
    .Y(_08604_));
 sky130_fd_sc_hd__a211o_4 _14745_ (.A1(_08346_),
    .A2(_08602_),
    .B1(_08444_),
    .C1(_08604_),
    .X(_00402_));
 sky130_fd_sc_hd__nor2_4 _14746_ (.A(\CPU_Xreg_value_a4[19][3] ),
    .B(_08532_),
    .Y(_08605_));
 sky130_fd_sc_hd__a211o_4 _14747_ (.A1(_08348_),
    .A2(_08535_),
    .B1(_08591_),
    .C1(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__inv_2 _14748_ (.A(_08606_),
    .Y(_00401_));
 sky130_fd_sc_hd__buf_2 _14749_ (.A(_08560_),
    .X(_08607_));
 sky130_fd_sc_hd__nor2_4 _14750_ (.A(\CPU_Xreg_value_a4[19][2] ),
    .B(_08532_),
    .Y(_08608_));
 sky130_fd_sc_hd__a211o_4 _14751_ (.A1(_08351_),
    .A2(_08535_),
    .B1(_08607_),
    .C1(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__inv_2 _14752_ (.A(_08609_),
    .Y(_00400_));
 sky130_fd_sc_hd__inv_2 _14753_ (.A(\CPU_Xreg_value_a4[19][1] ),
    .Y(_08610_));
 sky130_fd_sc_hd__nor2_4 _14754_ (.A(_08610_),
    .B(_08602_),
    .Y(_08611_));
 sky130_fd_sc_hd__a211o_4 _14755_ (.A1(_08181_),
    .A2(_08602_),
    .B1(_08444_),
    .C1(_08611_),
    .X(_00399_));
 sky130_fd_sc_hd__inv_2 _14756_ (.A(\CPU_Xreg_value_a4[19][0] ),
    .Y(_08612_));
 sky130_fd_sc_hd__nor2_4 _14757_ (.A(_08612_),
    .B(_08602_),
    .Y(_08613_));
 sky130_fd_sc_hd__a211o_4 _14758_ (.A1(_08270_),
    .A2(_08602_),
    .B1(_08444_),
    .C1(_08613_),
    .X(_00398_));
 sky130_fd_sc_hd__buf_2 _14759_ (.A(_06503_),
    .X(_08614_));
 sky130_fd_sc_hd__or2_4 _14760_ (.A(_07193_),
    .B(_08362_),
    .X(_08615_));
 sky130_fd_sc_hd__inv_2 _14761_ (.A(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__buf_2 _14762_ (.A(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__buf_2 _14763_ (.A(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__buf_2 _14764_ (.A(_08616_),
    .X(_08619_));
 sky130_fd_sc_hd__buf_2 _14765_ (.A(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_4 _14766_ (.A(\CPU_Xreg_value_a4[20][31] ),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__a211o_4 _14767_ (.A1(_08614_),
    .A2(_08618_),
    .B1(_08607_),
    .C1(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__inv_2 _14768_ (.A(_08622_),
    .Y(_00397_));
 sky130_fd_sc_hd__buf_2 _14769_ (.A(_06515_),
    .X(_08623_));
 sky130_fd_sc_hd__nor2_4 _14770_ (.A(\CPU_Xreg_value_a4[20][30] ),
    .B(_08620_),
    .Y(_08624_));
 sky130_fd_sc_hd__a211o_4 _14771_ (.A1(_08623_),
    .A2(_08618_),
    .B1(_08607_),
    .C1(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__inv_2 _14772_ (.A(_08625_),
    .Y(_00396_));
 sky130_fd_sc_hd__buf_2 _14773_ (.A(_06531_),
    .X(_08626_));
 sky130_fd_sc_hd__nor2_4 _14774_ (.A(\CPU_Xreg_value_a4[20][29] ),
    .B(_08620_),
    .Y(_08627_));
 sky130_fd_sc_hd__a211o_4 _14775_ (.A1(_08626_),
    .A2(_08618_),
    .B1(_08607_),
    .C1(_08627_),
    .X(_08628_));
 sky130_fd_sc_hd__inv_2 _14776_ (.A(_08628_),
    .Y(_00395_));
 sky130_fd_sc_hd__buf_2 _14777_ (.A(_06539_),
    .X(_08629_));
 sky130_fd_sc_hd__nor2_4 _14778_ (.A(\CPU_Xreg_value_a4[20][28] ),
    .B(_08620_),
    .Y(_08630_));
 sky130_fd_sc_hd__a211o_4 _14779_ (.A1(_08629_),
    .A2(_08618_),
    .B1(_08607_),
    .C1(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__inv_2 _14780_ (.A(_08631_),
    .Y(_00394_));
 sky130_fd_sc_hd__buf_2 _14781_ (.A(_06564_),
    .X(_08632_));
 sky130_fd_sc_hd__buf_2 _14782_ (.A(_08617_),
    .X(_08633_));
 sky130_fd_sc_hd__buf_2 _14783_ (.A(_08619_),
    .X(_08634_));
 sky130_fd_sc_hd__nor2_4 _14784_ (.A(\CPU_Xreg_value_a4[20][27] ),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__a211o_4 _14785_ (.A1(_08632_),
    .A2(_08633_),
    .B1(_08607_),
    .C1(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__inv_2 _14786_ (.A(_08636_),
    .Y(_00393_));
 sky130_fd_sc_hd__buf_2 _14787_ (.A(_06574_),
    .X(_08637_));
 sky130_fd_sc_hd__buf_2 _14788_ (.A(_08560_),
    .X(_08638_));
 sky130_fd_sc_hd__nor2_4 _14789_ (.A(\CPU_Xreg_value_a4[20][26] ),
    .B(_08634_),
    .Y(_08639_));
 sky130_fd_sc_hd__a211o_4 _14790_ (.A1(_08637_),
    .A2(_08633_),
    .B1(_08638_),
    .C1(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__inv_2 _14791_ (.A(_08640_),
    .Y(_00392_));
 sky130_fd_sc_hd__buf_2 _14792_ (.A(_06589_),
    .X(_08641_));
 sky130_fd_sc_hd__nor2_4 _14793_ (.A(\CPU_Xreg_value_a4[20][25] ),
    .B(_08634_),
    .Y(_08642_));
 sky130_fd_sc_hd__a211o_4 _14794_ (.A1(_08641_),
    .A2(_08633_),
    .B1(_08638_),
    .C1(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__inv_2 _14795_ (.A(_08643_),
    .Y(_00391_));
 sky130_fd_sc_hd__buf_2 _14796_ (.A(_06599_),
    .X(_08644_));
 sky130_fd_sc_hd__nor2_4 _14797_ (.A(\CPU_Xreg_value_a4[20][24] ),
    .B(_08634_),
    .Y(_08645_));
 sky130_fd_sc_hd__a211o_4 _14798_ (.A1(_08644_),
    .A2(_08633_),
    .B1(_08638_),
    .C1(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__inv_2 _14799_ (.A(_08646_),
    .Y(_00390_));
 sky130_fd_sc_hd__buf_2 _14800_ (.A(_06619_),
    .X(_08647_));
 sky130_fd_sc_hd__nor2_4 _14801_ (.A(\CPU_Xreg_value_a4[20][23] ),
    .B(_08634_),
    .Y(_08648_));
 sky130_fd_sc_hd__a211o_4 _14802_ (.A1(_08647_),
    .A2(_08633_),
    .B1(_08638_),
    .C1(_08648_),
    .X(_08649_));
 sky130_fd_sc_hd__inv_2 _14803_ (.A(_08649_),
    .Y(_00389_));
 sky130_fd_sc_hd__buf_2 _14804_ (.A(_06627_),
    .X(_08650_));
 sky130_fd_sc_hd__nor2_4 _14805_ (.A(\CPU_Xreg_value_a4[20][22] ),
    .B(_08634_),
    .Y(_08651_));
 sky130_fd_sc_hd__a211o_4 _14806_ (.A1(_08650_),
    .A2(_08633_),
    .B1(_08638_),
    .C1(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__inv_2 _14807_ (.A(_08652_),
    .Y(_00388_));
 sky130_fd_sc_hd__buf_2 _14808_ (.A(_06642_),
    .X(_08653_));
 sky130_fd_sc_hd__buf_2 _14809_ (.A(_08617_),
    .X(_08654_));
 sky130_fd_sc_hd__buf_2 _14810_ (.A(_08619_),
    .X(_08655_));
 sky130_fd_sc_hd__nor2_4 _14811_ (.A(\CPU_Xreg_value_a4[20][21] ),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__a211o_4 _14812_ (.A1(_08653_),
    .A2(_08654_),
    .B1(_08638_),
    .C1(_08656_),
    .X(_08657_));
 sky130_fd_sc_hd__inv_2 _14813_ (.A(_08657_),
    .Y(_00387_));
 sky130_fd_sc_hd__buf_2 _14814_ (.A(_06651_),
    .X(_08658_));
 sky130_fd_sc_hd__buf_2 _14815_ (.A(_08560_),
    .X(_08659_));
 sky130_fd_sc_hd__nor2_4 _14816_ (.A(\CPU_Xreg_value_a4[20][20] ),
    .B(_08655_),
    .Y(_08660_));
 sky130_fd_sc_hd__a211o_4 _14817_ (.A1(_08658_),
    .A2(_08654_),
    .B1(_08659_),
    .C1(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__inv_2 _14818_ (.A(_08661_),
    .Y(_00386_));
 sky130_fd_sc_hd__buf_2 _14819_ (.A(_06673_),
    .X(_08662_));
 sky130_fd_sc_hd__nor2_4 _14820_ (.A(\CPU_Xreg_value_a4[20][19] ),
    .B(_08655_),
    .Y(_08663_));
 sky130_fd_sc_hd__a211o_4 _14821_ (.A1(_08662_),
    .A2(_08654_),
    .B1(_08659_),
    .C1(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__inv_2 _14822_ (.A(_08664_),
    .Y(_00385_));
 sky130_fd_sc_hd__buf_2 _14823_ (.A(_06682_),
    .X(_08665_));
 sky130_fd_sc_hd__nor2_4 _14824_ (.A(\CPU_Xreg_value_a4[20][18] ),
    .B(_08655_),
    .Y(_08666_));
 sky130_fd_sc_hd__a211o_4 _14825_ (.A1(_08665_),
    .A2(_08654_),
    .B1(_08659_),
    .C1(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__inv_2 _14826_ (.A(_08667_),
    .Y(_00384_));
 sky130_fd_sc_hd__buf_2 _14827_ (.A(_06692_),
    .X(_08668_));
 sky130_fd_sc_hd__nor2_4 _14828_ (.A(\CPU_Xreg_value_a4[20][17] ),
    .B(_08655_),
    .Y(_08669_));
 sky130_fd_sc_hd__a211o_4 _14829_ (.A1(_08668_),
    .A2(_08654_),
    .B1(_08659_),
    .C1(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__inv_2 _14830_ (.A(_08670_),
    .Y(_00383_));
 sky130_fd_sc_hd__buf_2 _14831_ (.A(_06701_),
    .X(_08671_));
 sky130_fd_sc_hd__nor2_4 _14832_ (.A(\CPU_Xreg_value_a4[20][16] ),
    .B(_08655_),
    .Y(_08672_));
 sky130_fd_sc_hd__a211o_4 _14833_ (.A1(_08671_),
    .A2(_08654_),
    .B1(_08659_),
    .C1(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__inv_2 _14834_ (.A(_08673_),
    .Y(_00382_));
 sky130_fd_sc_hd__buf_2 _14835_ (.A(_06724_),
    .X(_08674_));
 sky130_fd_sc_hd__buf_2 _14836_ (.A(_08617_),
    .X(_08675_));
 sky130_fd_sc_hd__buf_2 _14837_ (.A(_08619_),
    .X(_08676_));
 sky130_fd_sc_hd__nor2_4 _14838_ (.A(\CPU_Xreg_value_a4[20][15] ),
    .B(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__a211o_4 _14839_ (.A1(_08674_),
    .A2(_08675_),
    .B1(_08659_),
    .C1(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__inv_2 _14840_ (.A(_08678_),
    .Y(_00381_));
 sky130_fd_sc_hd__buf_2 _14841_ (.A(_06733_),
    .X(_08679_));
 sky130_fd_sc_hd__buf_2 _14842_ (.A(_08462_),
    .X(_08680_));
 sky130_fd_sc_hd__buf_2 _14843_ (.A(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__nor2_4 _14844_ (.A(\CPU_Xreg_value_a4[20][14] ),
    .B(_08676_),
    .Y(_08682_));
 sky130_fd_sc_hd__a211o_4 _14845_ (.A1(_08679_),
    .A2(_08675_),
    .B1(_08681_),
    .C1(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__inv_2 _14846_ (.A(_08683_),
    .Y(_00380_));
 sky130_fd_sc_hd__buf_2 _14847_ (.A(_06743_),
    .X(_08684_));
 sky130_fd_sc_hd__nor2_4 _14848_ (.A(\CPU_Xreg_value_a4[20][13] ),
    .B(_08676_),
    .Y(_08685_));
 sky130_fd_sc_hd__a211o_4 _14849_ (.A1(_08684_),
    .A2(_08675_),
    .B1(_08681_),
    .C1(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__inv_2 _14850_ (.A(_08686_),
    .Y(_00379_));
 sky130_fd_sc_hd__buf_2 _14851_ (.A(_06752_),
    .X(_08687_));
 sky130_fd_sc_hd__nor2_4 _14852_ (.A(\CPU_Xreg_value_a4[20][12] ),
    .B(_08676_),
    .Y(_08688_));
 sky130_fd_sc_hd__a211o_4 _14853_ (.A1(_08687_),
    .A2(_08675_),
    .B1(_08681_),
    .C1(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__inv_2 _14854_ (.A(_08689_),
    .Y(_00378_));
 sky130_fd_sc_hd__buf_2 _14855_ (.A(_06770_),
    .X(_08690_));
 sky130_fd_sc_hd__nor2_4 _14856_ (.A(\CPU_Xreg_value_a4[20][11] ),
    .B(_08676_),
    .Y(_08691_));
 sky130_fd_sc_hd__a211o_4 _14857_ (.A1(_08690_),
    .A2(_08675_),
    .B1(_08681_),
    .C1(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__inv_2 _14858_ (.A(_08692_),
    .Y(_00377_));
 sky130_fd_sc_hd__buf_2 _14859_ (.A(_06778_),
    .X(_08693_));
 sky130_fd_sc_hd__nor2_4 _14860_ (.A(\CPU_Xreg_value_a4[20][10] ),
    .B(_08676_),
    .Y(_08694_));
 sky130_fd_sc_hd__a211o_4 _14861_ (.A1(_08693_),
    .A2(_08675_),
    .B1(_08681_),
    .C1(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__inv_2 _14862_ (.A(_08695_),
    .Y(_00376_));
 sky130_fd_sc_hd__buf_2 _14863_ (.A(_06791_),
    .X(_08696_));
 sky130_fd_sc_hd__buf_2 _14864_ (.A(_08619_),
    .X(_08697_));
 sky130_fd_sc_hd__buf_2 _14865_ (.A(_08619_),
    .X(_08698_));
 sky130_fd_sc_hd__nor2_4 _14866_ (.A(\CPU_Xreg_value_a4[20][9] ),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__a211o_4 _14867_ (.A1(_08696_),
    .A2(_08697_),
    .B1(_08681_),
    .C1(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__inv_2 _14868_ (.A(_08700_),
    .Y(_00375_));
 sky130_fd_sc_hd__buf_2 _14869_ (.A(_06799_),
    .X(_08701_));
 sky130_fd_sc_hd__buf_2 _14870_ (.A(_08680_),
    .X(_08702_));
 sky130_fd_sc_hd__nor2_4 _14871_ (.A(\CPU_Xreg_value_a4[20][8] ),
    .B(_08698_),
    .Y(_08703_));
 sky130_fd_sc_hd__a211o_4 _14872_ (.A1(_08701_),
    .A2(_08697_),
    .B1(_08702_),
    .C1(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__inv_2 _14873_ (.A(_08704_),
    .Y(_00374_));
 sky130_fd_sc_hd__buf_2 _14874_ (.A(_06820_),
    .X(_08705_));
 sky130_fd_sc_hd__nor2_4 _14875_ (.A(\CPU_Xreg_value_a4[20][7] ),
    .B(_08698_),
    .Y(_08706_));
 sky130_fd_sc_hd__a211o_4 _14876_ (.A1(_08705_),
    .A2(_08697_),
    .B1(_08702_),
    .C1(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__inv_2 _14877_ (.A(_08707_),
    .Y(_00373_));
 sky130_fd_sc_hd__buf_2 _14878_ (.A(_06828_),
    .X(_08708_));
 sky130_fd_sc_hd__nor2_4 _14879_ (.A(\CPU_Xreg_value_a4[20][6] ),
    .B(_08698_),
    .Y(_08709_));
 sky130_fd_sc_hd__a211o_4 _14880_ (.A1(_08708_),
    .A2(_08697_),
    .B1(_08702_),
    .C1(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__inv_2 _14881_ (.A(_08710_),
    .Y(_00372_));
 sky130_fd_sc_hd__buf_2 _14882_ (.A(_06837_),
    .X(_08711_));
 sky130_fd_sc_hd__nor2_4 _14883_ (.A(\CPU_Xreg_value_a4[20][5] ),
    .B(_08698_),
    .Y(_08712_));
 sky130_fd_sc_hd__a211o_4 _14884_ (.A1(_08711_),
    .A2(_08697_),
    .B1(_08702_),
    .C1(_08712_),
    .X(_08713_));
 sky130_fd_sc_hd__inv_2 _14885_ (.A(_08713_),
    .Y(_00371_));
 sky130_fd_sc_hd__buf_2 _14886_ (.A(_08065_),
    .X(_08714_));
 sky130_fd_sc_hd__and2_4 _14887_ (.A(\CPU_Xreg_value_a4[20][4] ),
    .B(_08615_),
    .X(_08715_));
 sky130_fd_sc_hd__a211o_4 _14888_ (.A1(_08346_),
    .A2(_08618_),
    .B1(_08714_),
    .C1(_08715_),
    .X(_00370_));
 sky130_fd_sc_hd__nor2_4 _14889_ (.A(\CPU_Xreg_value_a4[20][3] ),
    .B(_08698_),
    .Y(_08716_));
 sky130_fd_sc_hd__a211o_4 _14890_ (.A1(_08348_),
    .A2(_08697_),
    .B1(_08702_),
    .C1(_08716_),
    .X(_08717_));
 sky130_fd_sc_hd__inv_2 _14891_ (.A(_08717_),
    .Y(_00369_));
 sky130_fd_sc_hd__and2_4 _14892_ (.A(\CPU_Xreg_value_a4[20][2] ),
    .B(_08615_),
    .X(_08718_));
 sky130_fd_sc_hd__a211o_4 _14893_ (.A1(_08178_),
    .A2(_08618_),
    .B1(_08714_),
    .C1(_08718_),
    .X(_00368_));
 sky130_fd_sc_hd__nor2_4 _14894_ (.A(\CPU_Xreg_value_a4[20][1] ),
    .B(_08617_),
    .Y(_08719_));
 sky130_fd_sc_hd__a211o_4 _14895_ (.A1(_08354_),
    .A2(_08620_),
    .B1(_08702_),
    .C1(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__inv_2 _14896_ (.A(_08720_),
    .Y(_00367_));
 sky130_fd_sc_hd__buf_2 _14897_ (.A(_08680_),
    .X(_08721_));
 sky130_fd_sc_hd__nor2_4 _14898_ (.A(\CPU_Xreg_value_a4[20][0] ),
    .B(_08617_),
    .Y(_08722_));
 sky130_fd_sc_hd__a211o_4 _14899_ (.A1(_08184_),
    .A2(_08620_),
    .B1(_08721_),
    .C1(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__inv_2 _14900_ (.A(_08723_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_4 _14901_ (.A(_07282_),
    .B(_08363_),
    .Y(_08724_));
 sky130_fd_sc_hd__buf_2 _14902_ (.A(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__buf_2 _14903_ (.A(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__buf_2 _14904_ (.A(_08724_),
    .X(_08727_));
 sky130_fd_sc_hd__buf_2 _14905_ (.A(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__nor2_4 _14906_ (.A(\CPU_Xreg_value_a4[21][31] ),
    .B(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__a211o_4 _14907_ (.A1(_08614_),
    .A2(_08726_),
    .B1(_08721_),
    .C1(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__inv_2 _14908_ (.A(_08730_),
    .Y(_00365_));
 sky130_fd_sc_hd__buf_2 _14909_ (.A(_08727_),
    .X(_08731_));
 sky130_fd_sc_hd__nor2_4 _14910_ (.A(\CPU_Xreg_value_a4[21][30] ),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__a211o_4 _14911_ (.A1(_08623_),
    .A2(_08726_),
    .B1(_08721_),
    .C1(_08732_),
    .X(_08733_));
 sky130_fd_sc_hd__inv_2 _14912_ (.A(_08733_),
    .Y(_00364_));
 sky130_fd_sc_hd__nor2_4 _14913_ (.A(\CPU_Xreg_value_a4[21][29] ),
    .B(_08731_),
    .Y(_08734_));
 sky130_fd_sc_hd__a211o_4 _14914_ (.A1(_08626_),
    .A2(_08726_),
    .B1(_08721_),
    .C1(_08734_),
    .X(_08735_));
 sky130_fd_sc_hd__inv_2 _14915_ (.A(_08735_),
    .Y(_00363_));
 sky130_fd_sc_hd__nor2_4 _14916_ (.A(\CPU_Xreg_value_a4[21][28] ),
    .B(_08731_),
    .Y(_08736_));
 sky130_fd_sc_hd__a211o_4 _14917_ (.A1(_08629_),
    .A2(_08726_),
    .B1(_08721_),
    .C1(_08736_),
    .X(_08737_));
 sky130_fd_sc_hd__inv_2 _14918_ (.A(_08737_),
    .Y(_00362_));
 sky130_fd_sc_hd__nor2_4 _14919_ (.A(\CPU_Xreg_value_a4[21][27] ),
    .B(_08731_),
    .Y(_08738_));
 sky130_fd_sc_hd__a211o_4 _14920_ (.A1(_08632_),
    .A2(_08726_),
    .B1(_08721_),
    .C1(_08738_),
    .X(_08739_));
 sky130_fd_sc_hd__inv_2 _14921_ (.A(_08739_),
    .Y(_00361_));
 sky130_fd_sc_hd__buf_2 _14922_ (.A(_08680_),
    .X(_08740_));
 sky130_fd_sc_hd__nor2_4 _14923_ (.A(\CPU_Xreg_value_a4[21][26] ),
    .B(_08731_),
    .Y(_08741_));
 sky130_fd_sc_hd__a211o_4 _14924_ (.A1(_08637_),
    .A2(_08726_),
    .B1(_08740_),
    .C1(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__inv_2 _14925_ (.A(_08742_),
    .Y(_00360_));
 sky130_fd_sc_hd__buf_2 _14926_ (.A(_08727_),
    .X(_08743_));
 sky130_fd_sc_hd__nor2_4 _14927_ (.A(\CPU_Xreg_value_a4[21][25] ),
    .B(_08731_),
    .Y(_08744_));
 sky130_fd_sc_hd__a211o_4 _14928_ (.A1(_08641_),
    .A2(_08743_),
    .B1(_08740_),
    .C1(_08744_),
    .X(_08745_));
 sky130_fd_sc_hd__inv_2 _14929_ (.A(_08745_),
    .Y(_00359_));
 sky130_fd_sc_hd__buf_2 _14930_ (.A(_08727_),
    .X(_08746_));
 sky130_fd_sc_hd__nor2_4 _14931_ (.A(\CPU_Xreg_value_a4[21][24] ),
    .B(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__a211o_4 _14932_ (.A1(_08644_),
    .A2(_08743_),
    .B1(_08740_),
    .C1(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__inv_2 _14933_ (.A(_08748_),
    .Y(_00358_));
 sky130_fd_sc_hd__nor2_4 _14934_ (.A(\CPU_Xreg_value_a4[21][23] ),
    .B(_08746_),
    .Y(_08749_));
 sky130_fd_sc_hd__a211o_4 _14935_ (.A1(_08647_),
    .A2(_08743_),
    .B1(_08740_),
    .C1(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__inv_2 _14936_ (.A(_08750_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_4 _14937_ (.A(\CPU_Xreg_value_a4[21][22] ),
    .B(_08746_),
    .Y(_08751_));
 sky130_fd_sc_hd__a211o_4 _14938_ (.A1(_08650_),
    .A2(_08743_),
    .B1(_08740_),
    .C1(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__inv_2 _14939_ (.A(_08752_),
    .Y(_00356_));
 sky130_fd_sc_hd__nor2_4 _14940_ (.A(\CPU_Xreg_value_a4[21][21] ),
    .B(_08746_),
    .Y(_08753_));
 sky130_fd_sc_hd__a211o_4 _14941_ (.A1(_08653_),
    .A2(_08743_),
    .B1(_08740_),
    .C1(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__inv_2 _14942_ (.A(_08754_),
    .Y(_00355_));
 sky130_fd_sc_hd__buf_2 _14943_ (.A(_08680_),
    .X(_08755_));
 sky130_fd_sc_hd__nor2_4 _14944_ (.A(\CPU_Xreg_value_a4[21][20] ),
    .B(_08746_),
    .Y(_08756_));
 sky130_fd_sc_hd__a211o_4 _14945_ (.A1(_08658_),
    .A2(_08743_),
    .B1(_08755_),
    .C1(_08756_),
    .X(_08757_));
 sky130_fd_sc_hd__inv_2 _14946_ (.A(_08757_),
    .Y(_00354_));
 sky130_fd_sc_hd__buf_2 _14947_ (.A(_08727_),
    .X(_08758_));
 sky130_fd_sc_hd__nor2_4 _14948_ (.A(\CPU_Xreg_value_a4[21][19] ),
    .B(_08746_),
    .Y(_08759_));
 sky130_fd_sc_hd__a211o_4 _14949_ (.A1(_08662_),
    .A2(_08758_),
    .B1(_08755_),
    .C1(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__inv_2 _14950_ (.A(_08760_),
    .Y(_00353_));
 sky130_fd_sc_hd__buf_2 _14951_ (.A(_08724_),
    .X(_08761_));
 sky130_fd_sc_hd__nor2_4 _14952_ (.A(\CPU_Xreg_value_a4[21][18] ),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a211o_4 _14953_ (.A1(_08665_),
    .A2(_08758_),
    .B1(_08755_),
    .C1(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__inv_2 _14954_ (.A(_08763_),
    .Y(_00352_));
 sky130_fd_sc_hd__nor2_4 _14955_ (.A(\CPU_Xreg_value_a4[21][17] ),
    .B(_08761_),
    .Y(_08764_));
 sky130_fd_sc_hd__a211o_4 _14956_ (.A1(_08668_),
    .A2(_08758_),
    .B1(_08755_),
    .C1(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__inv_2 _14957_ (.A(_08765_),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_4 _14958_ (.A(\CPU_Xreg_value_a4[21][16] ),
    .B(_08761_),
    .Y(_08766_));
 sky130_fd_sc_hd__a211o_4 _14959_ (.A1(_08671_),
    .A2(_08758_),
    .B1(_08755_),
    .C1(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__inv_2 _14960_ (.A(_08767_),
    .Y(_00350_));
 sky130_fd_sc_hd__nor2_4 _14961_ (.A(\CPU_Xreg_value_a4[21][15] ),
    .B(_08761_),
    .Y(_08768_));
 sky130_fd_sc_hd__a211o_4 _14962_ (.A1(_08674_),
    .A2(_08758_),
    .B1(_08755_),
    .C1(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__inv_2 _14963_ (.A(_08769_),
    .Y(_00349_));
 sky130_fd_sc_hd__buf_2 _14964_ (.A(_08680_),
    .X(_08770_));
 sky130_fd_sc_hd__nor2_4 _14965_ (.A(\CPU_Xreg_value_a4[21][14] ),
    .B(_08761_),
    .Y(_08771_));
 sky130_fd_sc_hd__a211o_4 _14966_ (.A1(_08679_),
    .A2(_08758_),
    .B1(_08770_),
    .C1(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__inv_2 _14967_ (.A(_08772_),
    .Y(_00348_));
 sky130_fd_sc_hd__buf_2 _14968_ (.A(_08727_),
    .X(_08773_));
 sky130_fd_sc_hd__nor2_4 _14969_ (.A(\CPU_Xreg_value_a4[21][13] ),
    .B(_08761_),
    .Y(_08774_));
 sky130_fd_sc_hd__a211o_4 _14970_ (.A1(_08684_),
    .A2(_08773_),
    .B1(_08770_),
    .C1(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__inv_2 _14971_ (.A(_08775_),
    .Y(_00347_));
 sky130_fd_sc_hd__buf_2 _14972_ (.A(_08724_),
    .X(_08776_));
 sky130_fd_sc_hd__nor2_4 _14973_ (.A(\CPU_Xreg_value_a4[21][12] ),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__a211o_4 _14974_ (.A1(_08687_),
    .A2(_08773_),
    .B1(_08770_),
    .C1(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__inv_2 _14975_ (.A(_08778_),
    .Y(_00346_));
 sky130_fd_sc_hd__nor2_4 _14976_ (.A(\CPU_Xreg_value_a4[21][11] ),
    .B(_08776_),
    .Y(_08779_));
 sky130_fd_sc_hd__a211o_4 _14977_ (.A1(_08690_),
    .A2(_08773_),
    .B1(_08770_),
    .C1(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__inv_2 _14978_ (.A(_08780_),
    .Y(_00345_));
 sky130_fd_sc_hd__nor2_4 _14979_ (.A(\CPU_Xreg_value_a4[21][10] ),
    .B(_08776_),
    .Y(_08781_));
 sky130_fd_sc_hd__a211o_4 _14980_ (.A1(_08693_),
    .A2(_08773_),
    .B1(_08770_),
    .C1(_08781_),
    .X(_08782_));
 sky130_fd_sc_hd__inv_2 _14981_ (.A(_08782_),
    .Y(_00344_));
 sky130_fd_sc_hd__nor2_4 _14982_ (.A(\CPU_Xreg_value_a4[21][9] ),
    .B(_08776_),
    .Y(_08783_));
 sky130_fd_sc_hd__a211o_4 _14983_ (.A1(_08696_),
    .A2(_08773_),
    .B1(_08770_),
    .C1(_08783_),
    .X(_08784_));
 sky130_fd_sc_hd__inv_2 _14984_ (.A(_08784_),
    .Y(_00343_));
 sky130_fd_sc_hd__buf_2 _14985_ (.A(_08462_),
    .X(_08785_));
 sky130_fd_sc_hd__buf_2 _14986_ (.A(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__nor2_4 _14987_ (.A(\CPU_Xreg_value_a4[21][8] ),
    .B(_08776_),
    .Y(_08787_));
 sky130_fd_sc_hd__a211o_4 _14988_ (.A1(_08701_),
    .A2(_08773_),
    .B1(_08786_),
    .C1(_08787_),
    .X(_08788_));
 sky130_fd_sc_hd__inv_2 _14989_ (.A(_08788_),
    .Y(_00342_));
 sky130_fd_sc_hd__nor2_4 _14990_ (.A(\CPU_Xreg_value_a4[21][7] ),
    .B(_08776_),
    .Y(_08789_));
 sky130_fd_sc_hd__a211o_4 _14991_ (.A1(_08705_),
    .A2(_08728_),
    .B1(_08786_),
    .C1(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__inv_2 _14992_ (.A(_08790_),
    .Y(_00341_));
 sky130_fd_sc_hd__nor2_4 _14993_ (.A(\CPU_Xreg_value_a4[21][6] ),
    .B(_08725_),
    .Y(_08791_));
 sky130_fd_sc_hd__a211o_4 _14994_ (.A1(_08708_),
    .A2(_08728_),
    .B1(_08786_),
    .C1(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__inv_2 _14995_ (.A(_08792_),
    .Y(_00340_));
 sky130_fd_sc_hd__nor2_4 _14996_ (.A(\CPU_Xreg_value_a4[21][5] ),
    .B(_08725_),
    .Y(_08793_));
 sky130_fd_sc_hd__a211o_4 _14997_ (.A1(_08711_),
    .A2(_08728_),
    .B1(_08786_),
    .C1(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__inv_2 _14998_ (.A(_08794_),
    .Y(_00339_));
 sky130_fd_sc_hd__buf_2 _14999_ (.A(_08725_),
    .X(_08795_));
 sky130_fd_sc_hd__inv_2 _15000_ (.A(\CPU_Xreg_value_a4[21][4] ),
    .Y(_08796_));
 sky130_fd_sc_hd__nor2_4 _15001_ (.A(_08796_),
    .B(_08795_),
    .Y(_08797_));
 sky130_fd_sc_hd__a211o_4 _15002_ (.A1(_08346_),
    .A2(_08795_),
    .B1(_08714_),
    .C1(_08797_),
    .X(_00338_));
 sky130_fd_sc_hd__nor2_4 _15003_ (.A(\CPU_Xreg_value_a4[21][3] ),
    .B(_08725_),
    .Y(_08798_));
 sky130_fd_sc_hd__a211o_4 _15004_ (.A1(_08348_),
    .A2(_08728_),
    .B1(_08786_),
    .C1(_08798_),
    .X(_08799_));
 sky130_fd_sc_hd__inv_2 _15005_ (.A(_08799_),
    .Y(_00337_));
 sky130_fd_sc_hd__inv_2 _15006_ (.A(\CPU_Xreg_value_a4[21][2] ),
    .Y(_08800_));
 sky130_fd_sc_hd__nor2_4 _15007_ (.A(_08800_),
    .B(_08795_),
    .Y(_08801_));
 sky130_fd_sc_hd__a211o_4 _15008_ (.A1(_08178_),
    .A2(_08795_),
    .B1(_08714_),
    .C1(_08801_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_4 _15009_ (.A(\CPU_Xreg_value_a4[21][1] ),
    .B(_08725_),
    .Y(_08802_));
 sky130_fd_sc_hd__a211o_4 _15010_ (.A1(_08354_),
    .A2(_08728_),
    .B1(_08786_),
    .C1(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__inv_2 _15011_ (.A(_08803_),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _15012_ (.A(\CPU_Xreg_value_a4[21][0] ),
    .Y(_08804_));
 sky130_fd_sc_hd__nor2_4 _15013_ (.A(_08804_),
    .B(_08795_),
    .Y(_08805_));
 sky130_fd_sc_hd__a211o_4 _15014_ (.A1(_08270_),
    .A2(_08795_),
    .B1(_08714_),
    .C1(_08805_),
    .X(_00334_));
 sky130_fd_sc_hd__or2_4 _15015_ (.A(_07365_),
    .B(_08362_),
    .X(_08806_));
 sky130_fd_sc_hd__inv_2 _15016_ (.A(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__buf_2 _15017_ (.A(_08807_),
    .X(_08808_));
 sky130_fd_sc_hd__buf_2 _15018_ (.A(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__buf_2 _15019_ (.A(_08785_),
    .X(_08810_));
 sky130_fd_sc_hd__buf_2 _15020_ (.A(_08807_),
    .X(_08811_));
 sky130_fd_sc_hd__nor2_4 _15021_ (.A(\CPU_Xreg_value_a4[22][31] ),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__a211o_4 _15022_ (.A1(_08614_),
    .A2(_08809_),
    .B1(_08810_),
    .C1(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__inv_2 _15023_ (.A(_08813_),
    .Y(_00333_));
 sky130_fd_sc_hd__nor2_4 _15024_ (.A(\CPU_Xreg_value_a4[22][30] ),
    .B(_08811_),
    .Y(_08814_));
 sky130_fd_sc_hd__a211o_4 _15025_ (.A1(_08623_),
    .A2(_08809_),
    .B1(_08810_),
    .C1(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__inv_2 _15026_ (.A(_08815_),
    .Y(_00332_));
 sky130_fd_sc_hd__nor2_4 _15027_ (.A(\CPU_Xreg_value_a4[22][29] ),
    .B(_08811_),
    .Y(_08816_));
 sky130_fd_sc_hd__a211o_4 _15028_ (.A1(_08626_),
    .A2(_08809_),
    .B1(_08810_),
    .C1(_08816_),
    .X(_08817_));
 sky130_fd_sc_hd__inv_2 _15029_ (.A(_08817_),
    .Y(_00331_));
 sky130_fd_sc_hd__buf_2 _15030_ (.A(_08808_),
    .X(_08818_));
 sky130_fd_sc_hd__nor2_4 _15031_ (.A(\CPU_Xreg_value_a4[22][28] ),
    .B(_08811_),
    .Y(_08819_));
 sky130_fd_sc_hd__a211o_4 _15032_ (.A1(_08629_),
    .A2(_08818_),
    .B1(_08810_),
    .C1(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__inv_2 _15033_ (.A(_08820_),
    .Y(_00330_));
 sky130_fd_sc_hd__buf_2 _15034_ (.A(_08807_),
    .X(_08821_));
 sky130_fd_sc_hd__nor2_4 _15035_ (.A(\CPU_Xreg_value_a4[22][27] ),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__a211o_4 _15036_ (.A1(_08632_),
    .A2(_08818_),
    .B1(_08810_),
    .C1(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__inv_2 _15037_ (.A(_08823_),
    .Y(_00329_));
 sky130_fd_sc_hd__nor2_4 _15038_ (.A(\CPU_Xreg_value_a4[22][26] ),
    .B(_08821_),
    .Y(_08824_));
 sky130_fd_sc_hd__a211o_4 _15039_ (.A1(_08637_),
    .A2(_08818_),
    .B1(_08810_),
    .C1(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__inv_2 _15040_ (.A(_08825_),
    .Y(_00328_));
 sky130_fd_sc_hd__buf_2 _15041_ (.A(_08785_),
    .X(_08826_));
 sky130_fd_sc_hd__nor2_4 _15042_ (.A(\CPU_Xreg_value_a4[22][25] ),
    .B(_08821_),
    .Y(_08827_));
 sky130_fd_sc_hd__a211o_4 _15043_ (.A1(_08641_),
    .A2(_08818_),
    .B1(_08826_),
    .C1(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__inv_2 _15044_ (.A(_08828_),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_4 _15045_ (.A(\CPU_Xreg_value_a4[22][24] ),
    .B(_08821_),
    .Y(_08829_));
 sky130_fd_sc_hd__a211o_4 _15046_ (.A1(_08644_),
    .A2(_08818_),
    .B1(_08826_),
    .C1(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__inv_2 _15047_ (.A(_08830_),
    .Y(_00326_));
 sky130_fd_sc_hd__nor2_4 _15048_ (.A(\CPU_Xreg_value_a4[22][23] ),
    .B(_08821_),
    .Y(_08831_));
 sky130_fd_sc_hd__a211o_4 _15049_ (.A1(_08647_),
    .A2(_08818_),
    .B1(_08826_),
    .C1(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__inv_2 _15050_ (.A(_08832_),
    .Y(_00325_));
 sky130_fd_sc_hd__buf_2 _15051_ (.A(_08808_),
    .X(_08833_));
 sky130_fd_sc_hd__nor2_4 _15052_ (.A(\CPU_Xreg_value_a4[22][22] ),
    .B(_08821_),
    .Y(_08834_));
 sky130_fd_sc_hd__a211o_4 _15053_ (.A1(_08650_),
    .A2(_08833_),
    .B1(_08826_),
    .C1(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__inv_2 _15054_ (.A(_08835_),
    .Y(_00324_));
 sky130_fd_sc_hd__buf_2 _15055_ (.A(_08807_),
    .X(_08836_));
 sky130_fd_sc_hd__nor2_4 _15056_ (.A(\CPU_Xreg_value_a4[22][21] ),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__a211o_4 _15057_ (.A1(_08653_),
    .A2(_08833_),
    .B1(_08826_),
    .C1(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__inv_2 _15058_ (.A(_08838_),
    .Y(_00323_));
 sky130_fd_sc_hd__nor2_4 _15059_ (.A(\CPU_Xreg_value_a4[22][20] ),
    .B(_08836_),
    .Y(_08839_));
 sky130_fd_sc_hd__a211o_4 _15060_ (.A1(_08658_),
    .A2(_08833_),
    .B1(_08826_),
    .C1(_08839_),
    .X(_08840_));
 sky130_fd_sc_hd__inv_2 _15061_ (.A(_08840_),
    .Y(_00322_));
 sky130_fd_sc_hd__buf_2 _15062_ (.A(_08785_),
    .X(_08841_));
 sky130_fd_sc_hd__nor2_4 _15063_ (.A(\CPU_Xreg_value_a4[22][19] ),
    .B(_08836_),
    .Y(_08842_));
 sky130_fd_sc_hd__a211o_4 _15064_ (.A1(_08662_),
    .A2(_08833_),
    .B1(_08841_),
    .C1(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__inv_2 _15065_ (.A(_08843_),
    .Y(_00321_));
 sky130_fd_sc_hd__nor2_4 _15066_ (.A(\CPU_Xreg_value_a4[22][18] ),
    .B(_08836_),
    .Y(_08844_));
 sky130_fd_sc_hd__a211o_4 _15067_ (.A1(_08665_),
    .A2(_08833_),
    .B1(_08841_),
    .C1(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__inv_2 _15068_ (.A(_08845_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_4 _15069_ (.A(\CPU_Xreg_value_a4[22][17] ),
    .B(_08836_),
    .Y(_08846_));
 sky130_fd_sc_hd__a211o_4 _15070_ (.A1(_08668_),
    .A2(_08833_),
    .B1(_08841_),
    .C1(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__inv_2 _15071_ (.A(_08847_),
    .Y(_00319_));
 sky130_fd_sc_hd__buf_2 _15072_ (.A(_08808_),
    .X(_08848_));
 sky130_fd_sc_hd__nor2_4 _15073_ (.A(\CPU_Xreg_value_a4[22][16] ),
    .B(_08836_),
    .Y(_08849_));
 sky130_fd_sc_hd__a211o_4 _15074_ (.A1(_08671_),
    .A2(_08848_),
    .B1(_08841_),
    .C1(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__inv_2 _15075_ (.A(_08850_),
    .Y(_00318_));
 sky130_fd_sc_hd__buf_2 _15076_ (.A(_08807_),
    .X(_08851_));
 sky130_fd_sc_hd__nor2_4 _15077_ (.A(\CPU_Xreg_value_a4[22][15] ),
    .B(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__a211o_4 _15078_ (.A1(_08674_),
    .A2(_08848_),
    .B1(_08841_),
    .C1(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__inv_2 _15079_ (.A(_08853_),
    .Y(_00317_));
 sky130_fd_sc_hd__nor2_4 _15080_ (.A(\CPU_Xreg_value_a4[22][14] ),
    .B(_08851_),
    .Y(_08854_));
 sky130_fd_sc_hd__a211o_4 _15081_ (.A1(_08679_),
    .A2(_08848_),
    .B1(_08841_),
    .C1(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__inv_2 _15082_ (.A(_08855_),
    .Y(_00316_));
 sky130_fd_sc_hd__buf_2 _15083_ (.A(_08785_),
    .X(_08856_));
 sky130_fd_sc_hd__nor2_4 _15084_ (.A(\CPU_Xreg_value_a4[22][13] ),
    .B(_08851_),
    .Y(_08857_));
 sky130_fd_sc_hd__a211o_4 _15085_ (.A1(_08684_),
    .A2(_08848_),
    .B1(_08856_),
    .C1(_08857_),
    .X(_08858_));
 sky130_fd_sc_hd__inv_2 _15086_ (.A(_08858_),
    .Y(_00315_));
 sky130_fd_sc_hd__nor2_4 _15087_ (.A(\CPU_Xreg_value_a4[22][12] ),
    .B(_08851_),
    .Y(_08859_));
 sky130_fd_sc_hd__a211o_4 _15088_ (.A1(_08687_),
    .A2(_08848_),
    .B1(_08856_),
    .C1(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__inv_2 _15089_ (.A(_08860_),
    .Y(_00314_));
 sky130_fd_sc_hd__nor2_4 _15090_ (.A(\CPU_Xreg_value_a4[22][11] ),
    .B(_08851_),
    .Y(_08861_));
 sky130_fd_sc_hd__a211o_4 _15091_ (.A1(_08690_),
    .A2(_08848_),
    .B1(_08856_),
    .C1(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__inv_2 _15092_ (.A(_08862_),
    .Y(_00313_));
 sky130_fd_sc_hd__buf_2 _15093_ (.A(_08808_),
    .X(_08863_));
 sky130_fd_sc_hd__nor2_4 _15094_ (.A(\CPU_Xreg_value_a4[22][10] ),
    .B(_08851_),
    .Y(_08864_));
 sky130_fd_sc_hd__a211o_4 _15095_ (.A1(_08693_),
    .A2(_08863_),
    .B1(_08856_),
    .C1(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__inv_2 _15096_ (.A(_08865_),
    .Y(_00312_));
 sky130_fd_sc_hd__buf_2 _15097_ (.A(_08807_),
    .X(_08866_));
 sky130_fd_sc_hd__nor2_4 _15098_ (.A(\CPU_Xreg_value_a4[22][9] ),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__a211o_4 _15099_ (.A1(_08696_),
    .A2(_08863_),
    .B1(_08856_),
    .C1(_08867_),
    .X(_08868_));
 sky130_fd_sc_hd__inv_2 _15100_ (.A(_08868_),
    .Y(_00311_));
 sky130_fd_sc_hd__nor2_4 _15101_ (.A(\CPU_Xreg_value_a4[22][8] ),
    .B(_08866_),
    .Y(_08869_));
 sky130_fd_sc_hd__a211o_4 _15102_ (.A1(_08701_),
    .A2(_08863_),
    .B1(_08856_),
    .C1(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__inv_2 _15103_ (.A(_08870_),
    .Y(_00310_));
 sky130_fd_sc_hd__buf_2 _15104_ (.A(_08785_),
    .X(_08871_));
 sky130_fd_sc_hd__nor2_4 _15105_ (.A(\CPU_Xreg_value_a4[22][7] ),
    .B(_08866_),
    .Y(_08872_));
 sky130_fd_sc_hd__a211o_4 _15106_ (.A1(_08705_),
    .A2(_08863_),
    .B1(_08871_),
    .C1(_08872_),
    .X(_08873_));
 sky130_fd_sc_hd__inv_2 _15107_ (.A(_08873_),
    .Y(_00309_));
 sky130_fd_sc_hd__nor2_4 _15108_ (.A(\CPU_Xreg_value_a4[22][6] ),
    .B(_08866_),
    .Y(_08874_));
 sky130_fd_sc_hd__a211o_4 _15109_ (.A1(_08708_),
    .A2(_08863_),
    .B1(_08871_),
    .C1(_08874_),
    .X(_08875_));
 sky130_fd_sc_hd__inv_2 _15110_ (.A(_08875_),
    .Y(_00308_));
 sky130_fd_sc_hd__nor2_4 _15111_ (.A(\CPU_Xreg_value_a4[22][5] ),
    .B(_08866_),
    .Y(_08876_));
 sky130_fd_sc_hd__a211o_4 _15112_ (.A1(_08711_),
    .A2(_08863_),
    .B1(_08871_),
    .C1(_08876_),
    .X(_08877_));
 sky130_fd_sc_hd__inv_2 _15113_ (.A(_08877_),
    .Y(_00307_));
 sky130_fd_sc_hd__buf_2 _15114_ (.A(_08345_),
    .X(_08878_));
 sky130_fd_sc_hd__and2_4 _15115_ (.A(\CPU_Xreg_value_a4[22][4] ),
    .B(_08806_),
    .X(_08879_));
 sky130_fd_sc_hd__a211o_4 _15116_ (.A1(_08878_),
    .A2(_08809_),
    .B1(_08714_),
    .C1(_08879_),
    .X(_00306_));
 sky130_fd_sc_hd__nor2_4 _15117_ (.A(\CPU_Xreg_value_a4[22][3] ),
    .B(_08866_),
    .Y(_08880_));
 sky130_fd_sc_hd__a211o_4 _15118_ (.A1(_06852_),
    .A2(_08811_),
    .B1(_08871_),
    .C1(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__inv_2 _15119_ (.A(_08881_),
    .Y(_00305_));
 sky130_fd_sc_hd__buf_2 _15120_ (.A(_08065_),
    .X(_08882_));
 sky130_fd_sc_hd__and2_4 _15121_ (.A(\CPU_Xreg_value_a4[22][2] ),
    .B(_08806_),
    .X(_08883_));
 sky130_fd_sc_hd__a211o_4 _15122_ (.A1(_08178_),
    .A2(_08809_),
    .B1(_08882_),
    .C1(_08883_),
    .X(_00304_));
 sky130_fd_sc_hd__and2_4 _15123_ (.A(\CPU_Xreg_value_a4[22][1] ),
    .B(_08806_),
    .X(_08884_));
 sky130_fd_sc_hd__a211o_4 _15124_ (.A1(_08181_),
    .A2(_08809_),
    .B1(_08882_),
    .C1(_08884_),
    .X(_00303_));
 sky130_fd_sc_hd__nor2_4 _15125_ (.A(\CPU_Xreg_value_a4[22][0] ),
    .B(_08808_),
    .Y(_08885_));
 sky130_fd_sc_hd__a211o_4 _15126_ (.A1(_08184_),
    .A2(_08811_),
    .B1(_08871_),
    .C1(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__inv_2 _15127_ (.A(_08886_),
    .Y(_00302_));
 sky130_fd_sc_hd__or2_4 _15128_ (.A(_07450_),
    .B(_08361_),
    .X(_08887_));
 sky130_fd_sc_hd__inv_2 _15129_ (.A(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__buf_2 _15130_ (.A(_08888_),
    .X(_08889_));
 sky130_fd_sc_hd__buf_2 _15131_ (.A(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__buf_2 _15132_ (.A(_08889_),
    .X(_08891_));
 sky130_fd_sc_hd__nor2_4 _15133_ (.A(\CPU_Xreg_value_a4[23][31] ),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__a211o_4 _15134_ (.A1(_08614_),
    .A2(_08890_),
    .B1(_08871_),
    .C1(_08892_),
    .X(_08893_));
 sky130_fd_sc_hd__inv_2 _15135_ (.A(_08893_),
    .Y(_00301_));
 sky130_fd_sc_hd__buf_2 _15136_ (.A(_08462_),
    .X(_08894_));
 sky130_fd_sc_hd__buf_2 _15137_ (.A(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__nor2_4 _15138_ (.A(\CPU_Xreg_value_a4[23][30] ),
    .B(_08891_),
    .Y(_08896_));
 sky130_fd_sc_hd__a211o_4 _15139_ (.A1(_08623_),
    .A2(_08890_),
    .B1(_08895_),
    .C1(_08896_),
    .X(_08897_));
 sky130_fd_sc_hd__inv_2 _15140_ (.A(_08897_),
    .Y(_00300_));
 sky130_fd_sc_hd__buf_2 _15141_ (.A(_08889_),
    .X(_08898_));
 sky130_fd_sc_hd__nor2_4 _15142_ (.A(\CPU_Xreg_value_a4[23][29] ),
    .B(_08891_),
    .Y(_08899_));
 sky130_fd_sc_hd__a211o_4 _15143_ (.A1(_08626_),
    .A2(_08898_),
    .B1(_08895_),
    .C1(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__inv_2 _15144_ (.A(_08900_),
    .Y(_00299_));
 sky130_fd_sc_hd__nor2_4 _15145_ (.A(\CPU_Xreg_value_a4[23][28] ),
    .B(_08891_),
    .Y(_08901_));
 sky130_fd_sc_hd__a211o_4 _15146_ (.A1(_08629_),
    .A2(_08898_),
    .B1(_08895_),
    .C1(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__inv_2 _15147_ (.A(_08902_),
    .Y(_00298_));
 sky130_fd_sc_hd__buf_2 _15148_ (.A(_08888_),
    .X(_08903_));
 sky130_fd_sc_hd__nor2_4 _15149_ (.A(\CPU_Xreg_value_a4[23][27] ),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__a211o_4 _15150_ (.A1(_08632_),
    .A2(_08898_),
    .B1(_08895_),
    .C1(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__inv_2 _15151_ (.A(_08905_),
    .Y(_00297_));
 sky130_fd_sc_hd__nor2_4 _15152_ (.A(\CPU_Xreg_value_a4[23][26] ),
    .B(_08903_),
    .Y(_08906_));
 sky130_fd_sc_hd__a211o_4 _15153_ (.A1(_08637_),
    .A2(_08898_),
    .B1(_08895_),
    .C1(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__inv_2 _15154_ (.A(_08907_),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_4 _15155_ (.A(\CPU_Xreg_value_a4[23][25] ),
    .B(_08903_),
    .Y(_08908_));
 sky130_fd_sc_hd__a211o_4 _15156_ (.A1(_08641_),
    .A2(_08898_),
    .B1(_08895_),
    .C1(_08908_),
    .X(_08909_));
 sky130_fd_sc_hd__inv_2 _15157_ (.A(_08909_),
    .Y(_00295_));
 sky130_fd_sc_hd__buf_2 _15158_ (.A(_08894_),
    .X(_08910_));
 sky130_fd_sc_hd__nor2_4 _15159_ (.A(\CPU_Xreg_value_a4[23][24] ),
    .B(_08903_),
    .Y(_08911_));
 sky130_fd_sc_hd__a211o_4 _15160_ (.A1(_08644_),
    .A2(_08898_),
    .B1(_08910_),
    .C1(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__inv_2 _15161_ (.A(_08912_),
    .Y(_00294_));
 sky130_fd_sc_hd__buf_2 _15162_ (.A(_08889_),
    .X(_08913_));
 sky130_fd_sc_hd__nor2_4 _15163_ (.A(\CPU_Xreg_value_a4[23][23] ),
    .B(_08903_),
    .Y(_08914_));
 sky130_fd_sc_hd__a211o_4 _15164_ (.A1(_08647_),
    .A2(_08913_),
    .B1(_08910_),
    .C1(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__inv_2 _15165_ (.A(_08915_),
    .Y(_00293_));
 sky130_fd_sc_hd__nor2_4 _15166_ (.A(\CPU_Xreg_value_a4[23][22] ),
    .B(_08903_),
    .Y(_08916_));
 sky130_fd_sc_hd__a211o_4 _15167_ (.A1(_08650_),
    .A2(_08913_),
    .B1(_08910_),
    .C1(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__inv_2 _15168_ (.A(_08917_),
    .Y(_00292_));
 sky130_fd_sc_hd__buf_2 _15169_ (.A(_08888_),
    .X(_08918_));
 sky130_fd_sc_hd__nor2_4 _15170_ (.A(\CPU_Xreg_value_a4[23][21] ),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__a211o_4 _15171_ (.A1(_08653_),
    .A2(_08913_),
    .B1(_08910_),
    .C1(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__inv_2 _15172_ (.A(_08920_),
    .Y(_00291_));
 sky130_fd_sc_hd__nor2_4 _15173_ (.A(\CPU_Xreg_value_a4[23][20] ),
    .B(_08918_),
    .Y(_08921_));
 sky130_fd_sc_hd__a211o_4 _15174_ (.A1(_08658_),
    .A2(_08913_),
    .B1(_08910_),
    .C1(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__inv_2 _15175_ (.A(_08922_),
    .Y(_00290_));
 sky130_fd_sc_hd__nor2_4 _15176_ (.A(\CPU_Xreg_value_a4[23][19] ),
    .B(_08918_),
    .Y(_08923_));
 sky130_fd_sc_hd__a211o_4 _15177_ (.A1(_08662_),
    .A2(_08913_),
    .B1(_08910_),
    .C1(_08923_),
    .X(_08924_));
 sky130_fd_sc_hd__inv_2 _15178_ (.A(_08924_),
    .Y(_00289_));
 sky130_fd_sc_hd__buf_2 _15179_ (.A(_08894_),
    .X(_08925_));
 sky130_fd_sc_hd__nor2_4 _15180_ (.A(\CPU_Xreg_value_a4[23][18] ),
    .B(_08918_),
    .Y(_08926_));
 sky130_fd_sc_hd__a211o_4 _15181_ (.A1(_08665_),
    .A2(_08913_),
    .B1(_08925_),
    .C1(_08926_),
    .X(_08927_));
 sky130_fd_sc_hd__inv_2 _15182_ (.A(_08927_),
    .Y(_00288_));
 sky130_fd_sc_hd__buf_2 _15183_ (.A(_08889_),
    .X(_08928_));
 sky130_fd_sc_hd__nor2_4 _15184_ (.A(\CPU_Xreg_value_a4[23][17] ),
    .B(_08918_),
    .Y(_08929_));
 sky130_fd_sc_hd__a211o_4 _15185_ (.A1(_08668_),
    .A2(_08928_),
    .B1(_08925_),
    .C1(_08929_),
    .X(_08930_));
 sky130_fd_sc_hd__inv_2 _15186_ (.A(_08930_),
    .Y(_00287_));
 sky130_fd_sc_hd__nor2_4 _15187_ (.A(\CPU_Xreg_value_a4[23][16] ),
    .B(_08918_),
    .Y(_08931_));
 sky130_fd_sc_hd__a211o_4 _15188_ (.A1(_08671_),
    .A2(_08928_),
    .B1(_08925_),
    .C1(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__inv_2 _15189_ (.A(_08932_),
    .Y(_00286_));
 sky130_fd_sc_hd__buf_2 _15190_ (.A(_08888_),
    .X(_08933_));
 sky130_fd_sc_hd__nor2_4 _15191_ (.A(\CPU_Xreg_value_a4[23][15] ),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__a211o_4 _15192_ (.A1(_08674_),
    .A2(_08928_),
    .B1(_08925_),
    .C1(_08934_),
    .X(_08935_));
 sky130_fd_sc_hd__inv_2 _15193_ (.A(_08935_),
    .Y(_00285_));
 sky130_fd_sc_hd__nor2_4 _15194_ (.A(\CPU_Xreg_value_a4[23][14] ),
    .B(_08933_),
    .Y(_08936_));
 sky130_fd_sc_hd__a211o_4 _15195_ (.A1(_08679_),
    .A2(_08928_),
    .B1(_08925_),
    .C1(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__inv_2 _15196_ (.A(_08937_),
    .Y(_00284_));
 sky130_fd_sc_hd__nor2_4 _15197_ (.A(\CPU_Xreg_value_a4[23][13] ),
    .B(_08933_),
    .Y(_08938_));
 sky130_fd_sc_hd__a211o_4 _15198_ (.A1(_08684_),
    .A2(_08928_),
    .B1(_08925_),
    .C1(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__inv_2 _15199_ (.A(_08939_),
    .Y(_00283_));
 sky130_fd_sc_hd__buf_2 _15200_ (.A(_08894_),
    .X(_08940_));
 sky130_fd_sc_hd__nor2_4 _15201_ (.A(\CPU_Xreg_value_a4[23][12] ),
    .B(_08933_),
    .Y(_08941_));
 sky130_fd_sc_hd__a211o_4 _15202_ (.A1(_08687_),
    .A2(_08928_),
    .B1(_08940_),
    .C1(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__inv_2 _15203_ (.A(_08942_),
    .Y(_00282_));
 sky130_fd_sc_hd__buf_2 _15204_ (.A(_08889_),
    .X(_08943_));
 sky130_fd_sc_hd__nor2_4 _15205_ (.A(\CPU_Xreg_value_a4[23][11] ),
    .B(_08933_),
    .Y(_08944_));
 sky130_fd_sc_hd__a211o_4 _15206_ (.A1(_08690_),
    .A2(_08943_),
    .B1(_08940_),
    .C1(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__inv_2 _15207_ (.A(_08945_),
    .Y(_00281_));
 sky130_fd_sc_hd__nor2_4 _15208_ (.A(\CPU_Xreg_value_a4[23][10] ),
    .B(_08933_),
    .Y(_08946_));
 sky130_fd_sc_hd__a211o_4 _15209_ (.A1(_08693_),
    .A2(_08943_),
    .B1(_08940_),
    .C1(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__inv_2 _15210_ (.A(_08947_),
    .Y(_00280_));
 sky130_fd_sc_hd__buf_2 _15211_ (.A(_08888_),
    .X(_08948_));
 sky130_fd_sc_hd__nor2_4 _15212_ (.A(\CPU_Xreg_value_a4[23][9] ),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__a211o_4 _15213_ (.A1(_08696_),
    .A2(_08943_),
    .B1(_08940_),
    .C1(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__inv_2 _15214_ (.A(_08950_),
    .Y(_00279_));
 sky130_fd_sc_hd__nor2_4 _15215_ (.A(\CPU_Xreg_value_a4[23][8] ),
    .B(_08948_),
    .Y(_08951_));
 sky130_fd_sc_hd__a211o_4 _15216_ (.A1(_08701_),
    .A2(_08943_),
    .B1(_08940_),
    .C1(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__inv_2 _15217_ (.A(_08952_),
    .Y(_00278_));
 sky130_fd_sc_hd__nor2_4 _15218_ (.A(\CPU_Xreg_value_a4[23][7] ),
    .B(_08948_),
    .Y(_08953_));
 sky130_fd_sc_hd__a211o_4 _15219_ (.A1(_08705_),
    .A2(_08943_),
    .B1(_08940_),
    .C1(_08953_),
    .X(_08954_));
 sky130_fd_sc_hd__inv_2 _15220_ (.A(_08954_),
    .Y(_00277_));
 sky130_fd_sc_hd__buf_2 _15221_ (.A(_08894_),
    .X(_08955_));
 sky130_fd_sc_hd__nor2_4 _15222_ (.A(\CPU_Xreg_value_a4[23][6] ),
    .B(_08948_),
    .Y(_08956_));
 sky130_fd_sc_hd__a211o_4 _15223_ (.A1(_08708_),
    .A2(_08943_),
    .B1(_08955_),
    .C1(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__inv_2 _15224_ (.A(_08957_),
    .Y(_00276_));
 sky130_fd_sc_hd__nor2_4 _15225_ (.A(\CPU_Xreg_value_a4[23][5] ),
    .B(_08948_),
    .Y(_08958_));
 sky130_fd_sc_hd__a211o_4 _15226_ (.A1(_08711_),
    .A2(_08891_),
    .B1(_08955_),
    .C1(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__inv_2 _15227_ (.A(_08959_),
    .Y(_00275_));
 sky130_fd_sc_hd__and2_4 _15228_ (.A(\CPU_Xreg_value_a4[23][4] ),
    .B(_08887_),
    .X(_08960_));
 sky130_fd_sc_hd__a211o_4 _15229_ (.A1(_08878_),
    .A2(_08890_),
    .B1(_08882_),
    .C1(_08960_),
    .X(_00274_));
 sky130_fd_sc_hd__nor2_4 _15230_ (.A(\CPU_Xreg_value_a4[23][3] ),
    .B(_08948_),
    .Y(_08961_));
 sky130_fd_sc_hd__a211o_4 _15231_ (.A1(_06852_),
    .A2(_08891_),
    .B1(_08955_),
    .C1(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__inv_2 _15232_ (.A(_08962_),
    .Y(_00273_));
 sky130_fd_sc_hd__and2_4 _15233_ (.A(\CPU_Xreg_value_a4[23][2] ),
    .B(_08887_),
    .X(_08963_));
 sky130_fd_sc_hd__a211o_4 _15234_ (.A1(_08178_),
    .A2(_08890_),
    .B1(_08882_),
    .C1(_08963_),
    .X(_00272_));
 sky130_fd_sc_hd__and2_4 _15235_ (.A(\CPU_Xreg_value_a4[23][1] ),
    .B(_08887_),
    .X(_08964_));
 sky130_fd_sc_hd__a211o_4 _15236_ (.A1(_08181_),
    .A2(_08890_),
    .B1(_08882_),
    .C1(_08964_),
    .X(_00271_));
 sky130_fd_sc_hd__and2_4 _15237_ (.A(\CPU_Xreg_value_a4[23][0] ),
    .B(_08887_),
    .X(_08965_));
 sky130_fd_sc_hd__a211o_4 _15238_ (.A1(_08270_),
    .A2(_08890_),
    .B1(_08882_),
    .C1(_08965_),
    .X(_00270_));
 sky130_fd_sc_hd__or2_4 _15239_ (.A(_07538_),
    .B(_08362_),
    .X(_08966_));
 sky130_fd_sc_hd__inv_2 _15240_ (.A(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__buf_2 _15241_ (.A(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__buf_2 _15242_ (.A(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__buf_2 _15243_ (.A(_08967_),
    .X(_08970_));
 sky130_fd_sc_hd__buf_2 _15244_ (.A(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__nor2_4 _15245_ (.A(\CPU_Xreg_value_a4[24][31] ),
    .B(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__a211o_4 _15246_ (.A1(_08614_),
    .A2(_08969_),
    .B1(_08955_),
    .C1(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__inv_2 _15247_ (.A(_08973_),
    .Y(_00269_));
 sky130_fd_sc_hd__nor2_4 _15248_ (.A(\CPU_Xreg_value_a4[24][30] ),
    .B(_08971_),
    .Y(_08974_));
 sky130_fd_sc_hd__a211o_4 _15249_ (.A1(_08623_),
    .A2(_08969_),
    .B1(_08955_),
    .C1(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__inv_2 _15250_ (.A(_08975_),
    .Y(_00268_));
 sky130_fd_sc_hd__nor2_4 _15251_ (.A(\CPU_Xreg_value_a4[24][29] ),
    .B(_08971_),
    .Y(_08976_));
 sky130_fd_sc_hd__a211o_4 _15252_ (.A1(_08626_),
    .A2(_08969_),
    .B1(_08955_),
    .C1(_08976_),
    .X(_08977_));
 sky130_fd_sc_hd__inv_2 _15253_ (.A(_08977_),
    .Y(_00267_));
 sky130_fd_sc_hd__buf_2 _15254_ (.A(_08894_),
    .X(_08978_));
 sky130_fd_sc_hd__nor2_4 _15255_ (.A(\CPU_Xreg_value_a4[24][28] ),
    .B(_08971_),
    .Y(_08979_));
 sky130_fd_sc_hd__a211o_4 _15256_ (.A1(_08629_),
    .A2(_08969_),
    .B1(_08978_),
    .C1(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__inv_2 _15257_ (.A(_08980_),
    .Y(_00266_));
 sky130_fd_sc_hd__buf_2 _15258_ (.A(_08968_),
    .X(_08981_));
 sky130_fd_sc_hd__buf_2 _15259_ (.A(_08970_),
    .X(_08982_));
 sky130_fd_sc_hd__nor2_4 _15260_ (.A(\CPU_Xreg_value_a4[24][27] ),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__a211o_4 _15261_ (.A1(_08632_),
    .A2(_08981_),
    .B1(_08978_),
    .C1(_08983_),
    .X(_08984_));
 sky130_fd_sc_hd__inv_2 _15262_ (.A(_08984_),
    .Y(_00265_));
 sky130_fd_sc_hd__nor2_4 _15263_ (.A(\CPU_Xreg_value_a4[24][26] ),
    .B(_08982_),
    .Y(_08985_));
 sky130_fd_sc_hd__a211o_4 _15264_ (.A1(_08637_),
    .A2(_08981_),
    .B1(_08978_),
    .C1(_08985_),
    .X(_08986_));
 sky130_fd_sc_hd__inv_2 _15265_ (.A(_08986_),
    .Y(_00264_));
 sky130_fd_sc_hd__nor2_4 _15266_ (.A(\CPU_Xreg_value_a4[24][25] ),
    .B(_08982_),
    .Y(_08987_));
 sky130_fd_sc_hd__a211o_4 _15267_ (.A1(_08641_),
    .A2(_08981_),
    .B1(_08978_),
    .C1(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__inv_2 _15268_ (.A(_08988_),
    .Y(_00263_));
 sky130_fd_sc_hd__nor2_4 _15269_ (.A(\CPU_Xreg_value_a4[24][24] ),
    .B(_08982_),
    .Y(_08989_));
 sky130_fd_sc_hd__a211o_4 _15270_ (.A1(_08644_),
    .A2(_08981_),
    .B1(_08978_),
    .C1(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__inv_2 _15271_ (.A(_08990_),
    .Y(_00262_));
 sky130_fd_sc_hd__nor2_4 _15272_ (.A(\CPU_Xreg_value_a4[24][23] ),
    .B(_08982_),
    .Y(_08991_));
 sky130_fd_sc_hd__a211o_4 _15273_ (.A1(_08647_),
    .A2(_08981_),
    .B1(_08978_),
    .C1(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__inv_2 _15274_ (.A(_08992_),
    .Y(_00261_));
 sky130_fd_sc_hd__buf_2 _15275_ (.A(_08462_),
    .X(_08993_));
 sky130_fd_sc_hd__buf_2 _15276_ (.A(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__nor2_4 _15277_ (.A(\CPU_Xreg_value_a4[24][22] ),
    .B(_08982_),
    .Y(_08995_));
 sky130_fd_sc_hd__a211o_4 _15278_ (.A1(_08650_),
    .A2(_08981_),
    .B1(_08994_),
    .C1(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__inv_2 _15279_ (.A(_08996_),
    .Y(_00260_));
 sky130_fd_sc_hd__buf_2 _15280_ (.A(_08968_),
    .X(_08997_));
 sky130_fd_sc_hd__buf_2 _15281_ (.A(_08970_),
    .X(_08998_));
 sky130_fd_sc_hd__nor2_4 _15282_ (.A(\CPU_Xreg_value_a4[24][21] ),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__a211o_4 _15283_ (.A1(_08653_),
    .A2(_08997_),
    .B1(_08994_),
    .C1(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__inv_2 _15284_ (.A(_09000_),
    .Y(_00259_));
 sky130_fd_sc_hd__nor2_4 _15285_ (.A(\CPU_Xreg_value_a4[24][20] ),
    .B(_08998_),
    .Y(_09001_));
 sky130_fd_sc_hd__a211o_4 _15286_ (.A1(_08658_),
    .A2(_08997_),
    .B1(_08994_),
    .C1(_09001_),
    .X(_09002_));
 sky130_fd_sc_hd__inv_2 _15287_ (.A(_09002_),
    .Y(_00258_));
 sky130_fd_sc_hd__nor2_4 _15288_ (.A(\CPU_Xreg_value_a4[24][19] ),
    .B(_08998_),
    .Y(_09003_));
 sky130_fd_sc_hd__a211o_4 _15289_ (.A1(_08662_),
    .A2(_08997_),
    .B1(_08994_),
    .C1(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__inv_2 _15290_ (.A(_09004_),
    .Y(_00257_));
 sky130_fd_sc_hd__nor2_4 _15291_ (.A(\CPU_Xreg_value_a4[24][18] ),
    .B(_08998_),
    .Y(_09005_));
 sky130_fd_sc_hd__a211o_4 _15292_ (.A1(_08665_),
    .A2(_08997_),
    .B1(_08994_),
    .C1(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__inv_2 _15293_ (.A(_09006_),
    .Y(_00256_));
 sky130_fd_sc_hd__nor2_4 _15294_ (.A(\CPU_Xreg_value_a4[24][17] ),
    .B(_08998_),
    .Y(_09007_));
 sky130_fd_sc_hd__a211o_4 _15295_ (.A1(_08668_),
    .A2(_08997_),
    .B1(_08994_),
    .C1(_09007_),
    .X(_09008_));
 sky130_fd_sc_hd__inv_2 _15296_ (.A(_09008_),
    .Y(_00255_));
 sky130_fd_sc_hd__buf_2 _15297_ (.A(_08993_),
    .X(_09009_));
 sky130_fd_sc_hd__nor2_4 _15298_ (.A(\CPU_Xreg_value_a4[24][16] ),
    .B(_08998_),
    .Y(_09010_));
 sky130_fd_sc_hd__a211o_4 _15299_ (.A1(_08671_),
    .A2(_08997_),
    .B1(_09009_),
    .C1(_09010_),
    .X(_09011_));
 sky130_fd_sc_hd__inv_2 _15300_ (.A(_09011_),
    .Y(_00254_));
 sky130_fd_sc_hd__buf_2 _15301_ (.A(_08968_),
    .X(_09012_));
 sky130_fd_sc_hd__buf_2 _15302_ (.A(_08970_),
    .X(_09013_));
 sky130_fd_sc_hd__nor2_4 _15303_ (.A(\CPU_Xreg_value_a4[24][15] ),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__a211o_4 _15304_ (.A1(_08674_),
    .A2(_09012_),
    .B1(_09009_),
    .C1(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__inv_2 _15305_ (.A(_09015_),
    .Y(_00253_));
 sky130_fd_sc_hd__nor2_4 _15306_ (.A(\CPU_Xreg_value_a4[24][14] ),
    .B(_09013_),
    .Y(_09016_));
 sky130_fd_sc_hd__a211o_4 _15307_ (.A1(_08679_),
    .A2(_09012_),
    .B1(_09009_),
    .C1(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__inv_2 _15308_ (.A(_09017_),
    .Y(_00252_));
 sky130_fd_sc_hd__nor2_4 _15309_ (.A(\CPU_Xreg_value_a4[24][13] ),
    .B(_09013_),
    .Y(_09018_));
 sky130_fd_sc_hd__a211o_4 _15310_ (.A1(_08684_),
    .A2(_09012_),
    .B1(_09009_),
    .C1(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__inv_2 _15311_ (.A(_09019_),
    .Y(_00251_));
 sky130_fd_sc_hd__nor2_4 _15312_ (.A(\CPU_Xreg_value_a4[24][12] ),
    .B(_09013_),
    .Y(_09020_));
 sky130_fd_sc_hd__a211o_4 _15313_ (.A1(_08687_),
    .A2(_09012_),
    .B1(_09009_),
    .C1(_09020_),
    .X(_09021_));
 sky130_fd_sc_hd__inv_2 _15314_ (.A(_09021_),
    .Y(_00250_));
 sky130_fd_sc_hd__nor2_4 _15315_ (.A(\CPU_Xreg_value_a4[24][11] ),
    .B(_09013_),
    .Y(_09022_));
 sky130_fd_sc_hd__a211o_4 _15316_ (.A1(_08690_),
    .A2(_09012_),
    .B1(_09009_),
    .C1(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__inv_2 _15317_ (.A(_09023_),
    .Y(_00249_));
 sky130_fd_sc_hd__buf_2 _15318_ (.A(_08993_),
    .X(_09024_));
 sky130_fd_sc_hd__nor2_4 _15319_ (.A(\CPU_Xreg_value_a4[24][10] ),
    .B(_09013_),
    .Y(_09025_));
 sky130_fd_sc_hd__a211o_4 _15320_ (.A1(_08693_),
    .A2(_09012_),
    .B1(_09024_),
    .C1(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__inv_2 _15321_ (.A(_09026_),
    .Y(_00248_));
 sky130_fd_sc_hd__buf_2 _15322_ (.A(_08970_),
    .X(_09027_));
 sky130_fd_sc_hd__buf_2 _15323_ (.A(_08970_),
    .X(_09028_));
 sky130_fd_sc_hd__nor2_4 _15324_ (.A(\CPU_Xreg_value_a4[24][9] ),
    .B(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__a211o_4 _15325_ (.A1(_08696_),
    .A2(_09027_),
    .B1(_09024_),
    .C1(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__inv_2 _15326_ (.A(_09030_),
    .Y(_00247_));
 sky130_fd_sc_hd__nor2_4 _15327_ (.A(\CPU_Xreg_value_a4[24][8] ),
    .B(_09028_),
    .Y(_09031_));
 sky130_fd_sc_hd__a211o_4 _15328_ (.A1(_08701_),
    .A2(_09027_),
    .B1(_09024_),
    .C1(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__inv_2 _15329_ (.A(_09032_),
    .Y(_00246_));
 sky130_fd_sc_hd__nor2_4 _15330_ (.A(\CPU_Xreg_value_a4[24][7] ),
    .B(_09028_),
    .Y(_09033_));
 sky130_fd_sc_hd__a211o_4 _15331_ (.A1(_08705_),
    .A2(_09027_),
    .B1(_09024_),
    .C1(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__inv_2 _15332_ (.A(_09034_),
    .Y(_00245_));
 sky130_fd_sc_hd__nor2_4 _15333_ (.A(\CPU_Xreg_value_a4[24][6] ),
    .B(_09028_),
    .Y(_09035_));
 sky130_fd_sc_hd__a211o_4 _15334_ (.A1(_08708_),
    .A2(_09027_),
    .B1(_09024_),
    .C1(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__inv_2 _15335_ (.A(_09036_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_4 _15336_ (.A(\CPU_Xreg_value_a4[24][5] ),
    .B(_09028_),
    .Y(_09037_));
 sky130_fd_sc_hd__a211o_4 _15337_ (.A1(_08711_),
    .A2(_09027_),
    .B1(_09024_),
    .C1(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__inv_2 _15338_ (.A(_09038_),
    .Y(_00243_));
 sky130_fd_sc_hd__buf_2 _15339_ (.A(_08065_),
    .X(_09039_));
 sky130_fd_sc_hd__and2_4 _15340_ (.A(\CPU_Xreg_value_a4[24][4] ),
    .B(_08966_),
    .X(_09040_));
 sky130_fd_sc_hd__a211o_4 _15341_ (.A1(_08878_),
    .A2(_08969_),
    .B1(_09039_),
    .C1(_09040_),
    .X(_00242_));
 sky130_fd_sc_hd__and2_4 _15342_ (.A(\CPU_Xreg_value_a4[24][3] ),
    .B(_08966_),
    .X(_09041_));
 sky130_fd_sc_hd__a211o_4 _15343_ (.A1(_08174_),
    .A2(_08969_),
    .B1(_09039_),
    .C1(_09041_),
    .X(_00241_));
 sky130_fd_sc_hd__buf_2 _15344_ (.A(_08993_),
    .X(_09042_));
 sky130_fd_sc_hd__nor2_4 _15345_ (.A(\CPU_Xreg_value_a4[24][2] ),
    .B(_09028_),
    .Y(_09043_));
 sky130_fd_sc_hd__a211o_4 _15346_ (.A1(_08351_),
    .A2(_09027_),
    .B1(_09042_),
    .C1(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__inv_2 _15347_ (.A(_09044_),
    .Y(_00240_));
 sky130_fd_sc_hd__nor2_4 _15348_ (.A(\CPU_Xreg_value_a4[24][1] ),
    .B(_08968_),
    .Y(_09045_));
 sky130_fd_sc_hd__a211o_4 _15349_ (.A1(_08354_),
    .A2(_08971_),
    .B1(_09042_),
    .C1(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__inv_2 _15350_ (.A(_09046_),
    .Y(_00239_));
 sky130_fd_sc_hd__nor2_4 _15351_ (.A(\CPU_Xreg_value_a4[24][0] ),
    .B(_08968_),
    .Y(_09047_));
 sky130_fd_sc_hd__a211o_4 _15352_ (.A1(_08184_),
    .A2(_08971_),
    .B1(_09042_),
    .C1(_09047_),
    .X(_09048_));
 sky130_fd_sc_hd__inv_2 _15353_ (.A(_09048_),
    .Y(_00238_));
 sky130_fd_sc_hd__nor2_4 _15354_ (.A(_07651_),
    .B(_08363_),
    .Y(_09049_));
 sky130_fd_sc_hd__buf_2 _15355_ (.A(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__buf_2 _15356_ (.A(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__buf_2 _15357_ (.A(_09049_),
    .X(_09052_));
 sky130_fd_sc_hd__buf_2 _15358_ (.A(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__nor2_4 _15359_ (.A(\CPU_Xreg_value_a4[25][31] ),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__a211o_4 _15360_ (.A1(_08614_),
    .A2(_09051_),
    .B1(_09042_),
    .C1(_09054_),
    .X(_09055_));
 sky130_fd_sc_hd__inv_2 _15361_ (.A(_09055_),
    .Y(_00237_));
 sky130_fd_sc_hd__buf_2 _15362_ (.A(_09052_),
    .X(_09056_));
 sky130_fd_sc_hd__nor2_4 _15363_ (.A(\CPU_Xreg_value_a4[25][30] ),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__a211o_4 _15364_ (.A1(_08623_),
    .A2(_09051_),
    .B1(_09042_),
    .C1(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__inv_2 _15365_ (.A(_09058_),
    .Y(_00236_));
 sky130_fd_sc_hd__nor2_4 _15366_ (.A(\CPU_Xreg_value_a4[25][29] ),
    .B(_09056_),
    .Y(_09059_));
 sky130_fd_sc_hd__a211o_4 _15367_ (.A1(_08626_),
    .A2(_09051_),
    .B1(_09042_),
    .C1(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__inv_2 _15368_ (.A(_09060_),
    .Y(_00235_));
 sky130_fd_sc_hd__buf_2 _15369_ (.A(_08993_),
    .X(_09061_));
 sky130_fd_sc_hd__nor2_4 _15370_ (.A(\CPU_Xreg_value_a4[25][28] ),
    .B(_09056_),
    .Y(_09062_));
 sky130_fd_sc_hd__a211o_4 _15371_ (.A1(_08629_),
    .A2(_09051_),
    .B1(_09061_),
    .C1(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__inv_2 _15372_ (.A(_09063_),
    .Y(_00234_));
 sky130_fd_sc_hd__nor2_4 _15373_ (.A(\CPU_Xreg_value_a4[25][27] ),
    .B(_09056_),
    .Y(_09064_));
 sky130_fd_sc_hd__a211o_4 _15374_ (.A1(_08632_),
    .A2(_09051_),
    .B1(_09061_),
    .C1(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__inv_2 _15375_ (.A(_09065_),
    .Y(_00233_));
 sky130_fd_sc_hd__nor2_4 _15376_ (.A(\CPU_Xreg_value_a4[25][26] ),
    .B(_09056_),
    .Y(_09066_));
 sky130_fd_sc_hd__a211o_4 _15377_ (.A1(_08637_),
    .A2(_09051_),
    .B1(_09061_),
    .C1(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__inv_2 _15378_ (.A(_09067_),
    .Y(_00232_));
 sky130_fd_sc_hd__buf_2 _15379_ (.A(_09052_),
    .X(_09068_));
 sky130_fd_sc_hd__nor2_4 _15380_ (.A(\CPU_Xreg_value_a4[25][25] ),
    .B(_09056_),
    .Y(_09069_));
 sky130_fd_sc_hd__a211o_4 _15381_ (.A1(_08641_),
    .A2(_09068_),
    .B1(_09061_),
    .C1(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__inv_2 _15382_ (.A(_09070_),
    .Y(_00231_));
 sky130_fd_sc_hd__buf_2 _15383_ (.A(_09052_),
    .X(_09071_));
 sky130_fd_sc_hd__nor2_4 _15384_ (.A(\CPU_Xreg_value_a4[25][24] ),
    .B(_09071_),
    .Y(_09072_));
 sky130_fd_sc_hd__a211o_4 _15385_ (.A1(_08644_),
    .A2(_09068_),
    .B1(_09061_),
    .C1(_09072_),
    .X(_09073_));
 sky130_fd_sc_hd__inv_2 _15386_ (.A(_09073_),
    .Y(_00230_));
 sky130_fd_sc_hd__nor2_4 _15387_ (.A(\CPU_Xreg_value_a4[25][23] ),
    .B(_09071_),
    .Y(_09074_));
 sky130_fd_sc_hd__a211o_4 _15388_ (.A1(_08647_),
    .A2(_09068_),
    .B1(_09061_),
    .C1(_09074_),
    .X(_09075_));
 sky130_fd_sc_hd__inv_2 _15389_ (.A(_09075_),
    .Y(_00229_));
 sky130_fd_sc_hd__buf_2 _15390_ (.A(_08993_),
    .X(_09076_));
 sky130_fd_sc_hd__nor2_4 _15391_ (.A(\CPU_Xreg_value_a4[25][22] ),
    .B(_09071_),
    .Y(_09077_));
 sky130_fd_sc_hd__a211o_4 _15392_ (.A1(_08650_),
    .A2(_09068_),
    .B1(_09076_),
    .C1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__inv_2 _15393_ (.A(_09078_),
    .Y(_00228_));
 sky130_fd_sc_hd__nor2_4 _15394_ (.A(\CPU_Xreg_value_a4[25][21] ),
    .B(_09071_),
    .Y(_09079_));
 sky130_fd_sc_hd__a211o_4 _15395_ (.A1(_08653_),
    .A2(_09068_),
    .B1(_09076_),
    .C1(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__inv_2 _15396_ (.A(_09080_),
    .Y(_00227_));
 sky130_fd_sc_hd__nor2_4 _15397_ (.A(\CPU_Xreg_value_a4[25][20] ),
    .B(_09071_),
    .Y(_09081_));
 sky130_fd_sc_hd__a211o_4 _15398_ (.A1(_08658_),
    .A2(_09068_),
    .B1(_09076_),
    .C1(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__inv_2 _15399_ (.A(_09082_),
    .Y(_00226_));
 sky130_fd_sc_hd__buf_2 _15400_ (.A(_09052_),
    .X(_09083_));
 sky130_fd_sc_hd__nor2_4 _15401_ (.A(\CPU_Xreg_value_a4[25][19] ),
    .B(_09071_),
    .Y(_09084_));
 sky130_fd_sc_hd__a211o_4 _15402_ (.A1(_08662_),
    .A2(_09083_),
    .B1(_09076_),
    .C1(_09084_),
    .X(_09085_));
 sky130_fd_sc_hd__inv_2 _15403_ (.A(_09085_),
    .Y(_00225_));
 sky130_fd_sc_hd__buf_2 _15404_ (.A(_09049_),
    .X(_09086_));
 sky130_fd_sc_hd__nor2_4 _15405_ (.A(\CPU_Xreg_value_a4[25][18] ),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__a211o_4 _15406_ (.A1(_08665_),
    .A2(_09083_),
    .B1(_09076_),
    .C1(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__inv_2 _15407_ (.A(_09088_),
    .Y(_00224_));
 sky130_fd_sc_hd__nor2_4 _15408_ (.A(\CPU_Xreg_value_a4[25][17] ),
    .B(_09086_),
    .Y(_09089_));
 sky130_fd_sc_hd__a211o_4 _15409_ (.A1(_08668_),
    .A2(_09083_),
    .B1(_09076_),
    .C1(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__inv_2 _15410_ (.A(_09090_),
    .Y(_00223_));
 sky130_fd_sc_hd__buf_2 _15411_ (.A(_06100_),
    .X(_09091_));
 sky130_fd_sc_hd__buf_2 _15412_ (.A(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__nor2_4 _15413_ (.A(\CPU_Xreg_value_a4[25][16] ),
    .B(_09086_),
    .Y(_09093_));
 sky130_fd_sc_hd__a211o_4 _15414_ (.A1(_08671_),
    .A2(_09083_),
    .B1(_09092_),
    .C1(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__inv_2 _15415_ (.A(_09094_),
    .Y(_00222_));
 sky130_fd_sc_hd__nor2_4 _15416_ (.A(\CPU_Xreg_value_a4[25][15] ),
    .B(_09086_),
    .Y(_09095_));
 sky130_fd_sc_hd__a211o_4 _15417_ (.A1(_08674_),
    .A2(_09083_),
    .B1(_09092_),
    .C1(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__inv_2 _15418_ (.A(_09096_),
    .Y(_00221_));
 sky130_fd_sc_hd__nor2_4 _15419_ (.A(\CPU_Xreg_value_a4[25][14] ),
    .B(_09086_),
    .Y(_09097_));
 sky130_fd_sc_hd__a211o_4 _15420_ (.A1(_08679_),
    .A2(_09083_),
    .B1(_09092_),
    .C1(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__inv_2 _15421_ (.A(_09098_),
    .Y(_00220_));
 sky130_fd_sc_hd__buf_2 _15422_ (.A(_09052_),
    .X(_09099_));
 sky130_fd_sc_hd__nor2_4 _15423_ (.A(\CPU_Xreg_value_a4[25][13] ),
    .B(_09086_),
    .Y(_09100_));
 sky130_fd_sc_hd__a211o_4 _15424_ (.A1(_08684_),
    .A2(_09099_),
    .B1(_09092_),
    .C1(_09100_),
    .X(_09101_));
 sky130_fd_sc_hd__inv_2 _15425_ (.A(_09101_),
    .Y(_00219_));
 sky130_fd_sc_hd__buf_2 _15426_ (.A(_09049_),
    .X(_09102_));
 sky130_fd_sc_hd__nor2_4 _15427_ (.A(\CPU_Xreg_value_a4[25][12] ),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__a211o_4 _15428_ (.A1(_08687_),
    .A2(_09099_),
    .B1(_09092_),
    .C1(_09103_),
    .X(_09104_));
 sky130_fd_sc_hd__inv_2 _15429_ (.A(_09104_),
    .Y(_00218_));
 sky130_fd_sc_hd__nor2_4 _15430_ (.A(\CPU_Xreg_value_a4[25][11] ),
    .B(_09102_),
    .Y(_09105_));
 sky130_fd_sc_hd__a211o_4 _15431_ (.A1(_08690_),
    .A2(_09099_),
    .B1(_09092_),
    .C1(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__inv_2 _15432_ (.A(_09106_),
    .Y(_00217_));
 sky130_fd_sc_hd__buf_2 _15433_ (.A(_09091_),
    .X(_09107_));
 sky130_fd_sc_hd__nor2_4 _15434_ (.A(\CPU_Xreg_value_a4[25][10] ),
    .B(_09102_),
    .Y(_09108_));
 sky130_fd_sc_hd__a211o_4 _15435_ (.A1(_08693_),
    .A2(_09099_),
    .B1(_09107_),
    .C1(_09108_),
    .X(_09109_));
 sky130_fd_sc_hd__inv_2 _15436_ (.A(_09109_),
    .Y(_00216_));
 sky130_fd_sc_hd__nor2_4 _15437_ (.A(\CPU_Xreg_value_a4[25][9] ),
    .B(_09102_),
    .Y(_09110_));
 sky130_fd_sc_hd__a211o_4 _15438_ (.A1(_08696_),
    .A2(_09099_),
    .B1(_09107_),
    .C1(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__inv_2 _15439_ (.A(_09111_),
    .Y(_00215_));
 sky130_fd_sc_hd__nor2_4 _15440_ (.A(\CPU_Xreg_value_a4[25][8] ),
    .B(_09102_),
    .Y(_09112_));
 sky130_fd_sc_hd__a211o_4 _15441_ (.A1(_08701_),
    .A2(_09099_),
    .B1(_09107_),
    .C1(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__inv_2 _15442_ (.A(_09113_),
    .Y(_00214_));
 sky130_fd_sc_hd__nor2_4 _15443_ (.A(\CPU_Xreg_value_a4[25][7] ),
    .B(_09102_),
    .Y(_09114_));
 sky130_fd_sc_hd__a211o_4 _15444_ (.A1(_08705_),
    .A2(_09053_),
    .B1(_09107_),
    .C1(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__inv_2 _15445_ (.A(_09115_),
    .Y(_00213_));
 sky130_fd_sc_hd__nor2_4 _15446_ (.A(\CPU_Xreg_value_a4[25][6] ),
    .B(_09050_),
    .Y(_09116_));
 sky130_fd_sc_hd__a211o_4 _15447_ (.A1(_08708_),
    .A2(_09053_),
    .B1(_09107_),
    .C1(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__inv_2 _15448_ (.A(_09117_),
    .Y(_00212_));
 sky130_fd_sc_hd__nor2_4 _15449_ (.A(\CPU_Xreg_value_a4[25][5] ),
    .B(_09050_),
    .Y(_09118_));
 sky130_fd_sc_hd__a211o_4 _15450_ (.A1(_08711_),
    .A2(_09053_),
    .B1(_09107_),
    .C1(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__inv_2 _15451_ (.A(_09119_),
    .Y(_00211_));
 sky130_fd_sc_hd__buf_2 _15452_ (.A(_09050_),
    .X(_09120_));
 sky130_fd_sc_hd__inv_2 _15453_ (.A(\CPU_Xreg_value_a4[25][4] ),
    .Y(_09121_));
 sky130_fd_sc_hd__nor2_4 _15454_ (.A(_09121_),
    .B(_09120_),
    .Y(_09122_));
 sky130_fd_sc_hd__a211o_4 _15455_ (.A1(_08878_),
    .A2(_09120_),
    .B1(_09039_),
    .C1(_09122_),
    .X(_00210_));
 sky130_fd_sc_hd__inv_2 _15456_ (.A(\CPU_Xreg_value_a4[25][3] ),
    .Y(_09123_));
 sky130_fd_sc_hd__nor2_4 _15457_ (.A(_09123_),
    .B(_09120_),
    .Y(_09124_));
 sky130_fd_sc_hd__a211o_4 _15458_ (.A1(_08174_),
    .A2(_09120_),
    .B1(_09039_),
    .C1(_09124_),
    .X(_00209_));
 sky130_fd_sc_hd__buf_2 _15459_ (.A(_09091_),
    .X(_09125_));
 sky130_fd_sc_hd__nor2_4 _15460_ (.A(\CPU_Xreg_value_a4[25][2] ),
    .B(_09050_),
    .Y(_09126_));
 sky130_fd_sc_hd__a211o_4 _15461_ (.A1(_08351_),
    .A2(_09053_),
    .B1(_09125_),
    .C1(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__inv_2 _15462_ (.A(_09127_),
    .Y(_00208_));
 sky130_fd_sc_hd__nor2_4 _15463_ (.A(\CPU_Xreg_value_a4[25][1] ),
    .B(_09050_),
    .Y(_09128_));
 sky130_fd_sc_hd__a211o_4 _15464_ (.A1(_08354_),
    .A2(_09053_),
    .B1(_09125_),
    .C1(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__inv_2 _15465_ (.A(_09129_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _15466_ (.A(\CPU_Xreg_value_a4[25][0] ),
    .Y(_09130_));
 sky130_fd_sc_hd__nor2_4 _15467_ (.A(_09130_),
    .B(_09120_),
    .Y(_09131_));
 sky130_fd_sc_hd__a211o_4 _15468_ (.A1(_08270_),
    .A2(_09120_),
    .B1(_09039_),
    .C1(_09131_),
    .X(_00206_));
 sky130_fd_sc_hd__buf_2 _15469_ (.A(_06503_),
    .X(_09132_));
 sky130_fd_sc_hd__nor2_4 _15470_ (.A(_07735_),
    .B(_08363_),
    .Y(_09133_));
 sky130_fd_sc_hd__buf_2 _15471_ (.A(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__buf_2 _15472_ (.A(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__buf_2 _15473_ (.A(_09133_),
    .X(_09136_));
 sky130_fd_sc_hd__buf_2 _15474_ (.A(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__nor2_4 _15475_ (.A(\CPU_Xreg_value_a4[26][31] ),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__a211o_4 _15476_ (.A1(_09132_),
    .A2(_09135_),
    .B1(_09125_),
    .C1(_09138_),
    .X(_09139_));
 sky130_fd_sc_hd__inv_2 _15477_ (.A(_09139_),
    .Y(_00205_));
 sky130_fd_sc_hd__buf_2 _15478_ (.A(_06515_),
    .X(_09140_));
 sky130_fd_sc_hd__buf_2 _15479_ (.A(_09136_),
    .X(_09141_));
 sky130_fd_sc_hd__nor2_4 _15480_ (.A(\CPU_Xreg_value_a4[26][30] ),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__a211o_4 _15481_ (.A1(_09140_),
    .A2(_09135_),
    .B1(_09125_),
    .C1(_09142_),
    .X(_09143_));
 sky130_fd_sc_hd__inv_2 _15482_ (.A(_09143_),
    .Y(_00204_));
 sky130_fd_sc_hd__buf_2 _15483_ (.A(_06531_),
    .X(_09144_));
 sky130_fd_sc_hd__nor2_4 _15484_ (.A(\CPU_Xreg_value_a4[26][29] ),
    .B(_09141_),
    .Y(_09145_));
 sky130_fd_sc_hd__a211o_4 _15485_ (.A1(_09144_),
    .A2(_09135_),
    .B1(_09125_),
    .C1(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__inv_2 _15486_ (.A(_09146_),
    .Y(_00203_));
 sky130_fd_sc_hd__buf_2 _15487_ (.A(_06539_),
    .X(_09147_));
 sky130_fd_sc_hd__nor2_4 _15488_ (.A(\CPU_Xreg_value_a4[26][28] ),
    .B(_09141_),
    .Y(_09148_));
 sky130_fd_sc_hd__a211o_4 _15489_ (.A1(_09147_),
    .A2(_09135_),
    .B1(_09125_),
    .C1(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__inv_2 _15490_ (.A(_09149_),
    .Y(_00202_));
 sky130_fd_sc_hd__buf_2 _15491_ (.A(_06564_),
    .X(_09150_));
 sky130_fd_sc_hd__buf_2 _15492_ (.A(_09091_),
    .X(_09151_));
 sky130_fd_sc_hd__nor2_4 _15493_ (.A(\CPU_Xreg_value_a4[26][27] ),
    .B(_09141_),
    .Y(_09152_));
 sky130_fd_sc_hd__a211o_4 _15494_ (.A1(_09150_),
    .A2(_09135_),
    .B1(_09151_),
    .C1(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__inv_2 _15495_ (.A(_09153_),
    .Y(_00201_));
 sky130_fd_sc_hd__buf_2 _15496_ (.A(_06574_),
    .X(_09154_));
 sky130_fd_sc_hd__nor2_4 _15497_ (.A(\CPU_Xreg_value_a4[26][26] ),
    .B(_09141_),
    .Y(_09155_));
 sky130_fd_sc_hd__a211o_4 _15498_ (.A1(_09154_),
    .A2(_09135_),
    .B1(_09151_),
    .C1(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__inv_2 _15499_ (.A(_09156_),
    .Y(_00200_));
 sky130_fd_sc_hd__buf_2 _15500_ (.A(_06589_),
    .X(_09157_));
 sky130_fd_sc_hd__buf_2 _15501_ (.A(_09136_),
    .X(_09158_));
 sky130_fd_sc_hd__nor2_4 _15502_ (.A(\CPU_Xreg_value_a4[26][25] ),
    .B(_09141_),
    .Y(_09159_));
 sky130_fd_sc_hd__a211o_4 _15503_ (.A1(_09157_),
    .A2(_09158_),
    .B1(_09151_),
    .C1(_09159_),
    .X(_09160_));
 sky130_fd_sc_hd__inv_2 _15504_ (.A(_09160_),
    .Y(_00199_));
 sky130_fd_sc_hd__buf_2 _15505_ (.A(_06599_),
    .X(_09161_));
 sky130_fd_sc_hd__buf_2 _15506_ (.A(_09136_),
    .X(_09162_));
 sky130_fd_sc_hd__nor2_4 _15507_ (.A(\CPU_Xreg_value_a4[26][24] ),
    .B(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__a211o_4 _15508_ (.A1(_09161_),
    .A2(_09158_),
    .B1(_09151_),
    .C1(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__inv_2 _15509_ (.A(_09164_),
    .Y(_00198_));
 sky130_fd_sc_hd__buf_2 _15510_ (.A(_06619_),
    .X(_09165_));
 sky130_fd_sc_hd__nor2_4 _15511_ (.A(\CPU_Xreg_value_a4[26][23] ),
    .B(_09162_),
    .Y(_09166_));
 sky130_fd_sc_hd__a211o_4 _15512_ (.A1(_09165_),
    .A2(_09158_),
    .B1(_09151_),
    .C1(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__inv_2 _15513_ (.A(_09167_),
    .Y(_00197_));
 sky130_fd_sc_hd__buf_2 _15514_ (.A(_06627_),
    .X(_09168_));
 sky130_fd_sc_hd__nor2_4 _15515_ (.A(\CPU_Xreg_value_a4[26][22] ),
    .B(_09162_),
    .Y(_09169_));
 sky130_fd_sc_hd__a211o_4 _15516_ (.A1(_09168_),
    .A2(_09158_),
    .B1(_09151_),
    .C1(_09169_),
    .X(_09170_));
 sky130_fd_sc_hd__inv_2 _15517_ (.A(_09170_),
    .Y(_00196_));
 sky130_fd_sc_hd__buf_2 _15518_ (.A(_06642_),
    .X(_09171_));
 sky130_fd_sc_hd__buf_2 _15519_ (.A(_09091_),
    .X(_09172_));
 sky130_fd_sc_hd__nor2_4 _15520_ (.A(\CPU_Xreg_value_a4[26][21] ),
    .B(_09162_),
    .Y(_09173_));
 sky130_fd_sc_hd__a211o_4 _15521_ (.A1(_09171_),
    .A2(_09158_),
    .B1(_09172_),
    .C1(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__inv_2 _15522_ (.A(_09174_),
    .Y(_00195_));
 sky130_fd_sc_hd__buf_2 _15523_ (.A(_06651_),
    .X(_09175_));
 sky130_fd_sc_hd__nor2_4 _15524_ (.A(\CPU_Xreg_value_a4[26][20] ),
    .B(_09162_),
    .Y(_09176_));
 sky130_fd_sc_hd__a211o_4 _15525_ (.A1(_09175_),
    .A2(_09158_),
    .B1(_09172_),
    .C1(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__inv_2 _15526_ (.A(_09177_),
    .Y(_00194_));
 sky130_fd_sc_hd__buf_2 _15527_ (.A(_06673_),
    .X(_09178_));
 sky130_fd_sc_hd__buf_2 _15528_ (.A(_09136_),
    .X(_09179_));
 sky130_fd_sc_hd__nor2_4 _15529_ (.A(\CPU_Xreg_value_a4[26][19] ),
    .B(_09162_),
    .Y(_09180_));
 sky130_fd_sc_hd__a211o_4 _15530_ (.A1(_09178_),
    .A2(_09179_),
    .B1(_09172_),
    .C1(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__inv_2 _15531_ (.A(_09181_),
    .Y(_00193_));
 sky130_fd_sc_hd__buf_2 _15532_ (.A(_06682_),
    .X(_09182_));
 sky130_fd_sc_hd__buf_2 _15533_ (.A(_09133_),
    .X(_09183_));
 sky130_fd_sc_hd__nor2_4 _15534_ (.A(\CPU_Xreg_value_a4[26][18] ),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__a211o_4 _15535_ (.A1(_09182_),
    .A2(_09179_),
    .B1(_09172_),
    .C1(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__inv_2 _15536_ (.A(_09185_),
    .Y(_00192_));
 sky130_fd_sc_hd__buf_2 _15537_ (.A(_06692_),
    .X(_09186_));
 sky130_fd_sc_hd__nor2_4 _15538_ (.A(\CPU_Xreg_value_a4[26][17] ),
    .B(_09183_),
    .Y(_09187_));
 sky130_fd_sc_hd__a211o_4 _15539_ (.A1(_09186_),
    .A2(_09179_),
    .B1(_09172_),
    .C1(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__inv_2 _15540_ (.A(_09188_),
    .Y(_00191_));
 sky130_fd_sc_hd__buf_2 _15541_ (.A(_06701_),
    .X(_09189_));
 sky130_fd_sc_hd__nor2_4 _15542_ (.A(\CPU_Xreg_value_a4[26][16] ),
    .B(_09183_),
    .Y(_09190_));
 sky130_fd_sc_hd__a211o_4 _15543_ (.A1(_09189_),
    .A2(_09179_),
    .B1(_09172_),
    .C1(_09190_),
    .X(_09191_));
 sky130_fd_sc_hd__inv_2 _15544_ (.A(_09191_),
    .Y(_00190_));
 sky130_fd_sc_hd__buf_2 _15545_ (.A(_06724_),
    .X(_09192_));
 sky130_fd_sc_hd__buf_2 _15546_ (.A(_09091_),
    .X(_09193_));
 sky130_fd_sc_hd__nor2_4 _15547_ (.A(\CPU_Xreg_value_a4[26][15] ),
    .B(_09183_),
    .Y(_09194_));
 sky130_fd_sc_hd__a211o_4 _15548_ (.A1(_09192_),
    .A2(_09179_),
    .B1(_09193_),
    .C1(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__inv_2 _15549_ (.A(_09195_),
    .Y(_00189_));
 sky130_fd_sc_hd__buf_2 _15550_ (.A(_06733_),
    .X(_09196_));
 sky130_fd_sc_hd__nor2_4 _15551_ (.A(\CPU_Xreg_value_a4[26][14] ),
    .B(_09183_),
    .Y(_09197_));
 sky130_fd_sc_hd__a211o_4 _15552_ (.A1(_09196_),
    .A2(_09179_),
    .B1(_09193_),
    .C1(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__inv_2 _15553_ (.A(_09198_),
    .Y(_00188_));
 sky130_fd_sc_hd__buf_2 _15554_ (.A(_06743_),
    .X(_09199_));
 sky130_fd_sc_hd__buf_2 _15555_ (.A(_09136_),
    .X(_09200_));
 sky130_fd_sc_hd__nor2_4 _15556_ (.A(\CPU_Xreg_value_a4[26][13] ),
    .B(_09183_),
    .Y(_09201_));
 sky130_fd_sc_hd__a211o_4 _15557_ (.A1(_09199_),
    .A2(_09200_),
    .B1(_09193_),
    .C1(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__inv_2 _15558_ (.A(_09202_),
    .Y(_00187_));
 sky130_fd_sc_hd__buf_2 _15559_ (.A(_06752_),
    .X(_09203_));
 sky130_fd_sc_hd__buf_2 _15560_ (.A(_09133_),
    .X(_09204_));
 sky130_fd_sc_hd__nor2_4 _15561_ (.A(\CPU_Xreg_value_a4[26][12] ),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__a211o_4 _15562_ (.A1(_09203_),
    .A2(_09200_),
    .B1(_09193_),
    .C1(_09205_),
    .X(_09206_));
 sky130_fd_sc_hd__inv_2 _15563_ (.A(_09206_),
    .Y(_00186_));
 sky130_fd_sc_hd__buf_2 _15564_ (.A(_06770_),
    .X(_09207_));
 sky130_fd_sc_hd__nor2_4 _15565_ (.A(\CPU_Xreg_value_a4[26][11] ),
    .B(_09204_),
    .Y(_09208_));
 sky130_fd_sc_hd__a211o_4 _15566_ (.A1(_09207_),
    .A2(_09200_),
    .B1(_09193_),
    .C1(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__inv_2 _15567_ (.A(_09209_),
    .Y(_00185_));
 sky130_fd_sc_hd__buf_2 _15568_ (.A(_06778_),
    .X(_09210_));
 sky130_fd_sc_hd__nor2_4 _15569_ (.A(\CPU_Xreg_value_a4[26][10] ),
    .B(_09204_),
    .Y(_09211_));
 sky130_fd_sc_hd__a211o_4 _15570_ (.A1(_09210_),
    .A2(_09200_),
    .B1(_09193_),
    .C1(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__inv_2 _15571_ (.A(_09212_),
    .Y(_00184_));
 sky130_fd_sc_hd__buf_2 _15572_ (.A(_06791_),
    .X(_09213_));
 sky130_fd_sc_hd__buf_2 _15573_ (.A(_06100_),
    .X(_09214_));
 sky130_fd_sc_hd__buf_2 _15574_ (.A(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__nor2_4 _15575_ (.A(\CPU_Xreg_value_a4[26][9] ),
    .B(_09204_),
    .Y(_09216_));
 sky130_fd_sc_hd__a211o_4 _15576_ (.A1(_09213_),
    .A2(_09200_),
    .B1(_09215_),
    .C1(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__inv_2 _15577_ (.A(_09217_),
    .Y(_00183_));
 sky130_fd_sc_hd__buf_2 _15578_ (.A(_06799_),
    .X(_09218_));
 sky130_fd_sc_hd__nor2_4 _15579_ (.A(\CPU_Xreg_value_a4[26][8] ),
    .B(_09204_),
    .Y(_09219_));
 sky130_fd_sc_hd__a211o_4 _15580_ (.A1(_09218_),
    .A2(_09200_),
    .B1(_09215_),
    .C1(_09219_),
    .X(_09220_));
 sky130_fd_sc_hd__inv_2 _15581_ (.A(_09220_),
    .Y(_00182_));
 sky130_fd_sc_hd__buf_2 _15582_ (.A(_06820_),
    .X(_09221_));
 sky130_fd_sc_hd__nor2_4 _15583_ (.A(\CPU_Xreg_value_a4[26][7] ),
    .B(_09204_),
    .Y(_09222_));
 sky130_fd_sc_hd__a211o_4 _15584_ (.A1(_09221_),
    .A2(_09137_),
    .B1(_09215_),
    .C1(_09222_),
    .X(_09223_));
 sky130_fd_sc_hd__inv_2 _15585_ (.A(_09223_),
    .Y(_00181_));
 sky130_fd_sc_hd__buf_2 _15586_ (.A(_06828_),
    .X(_09224_));
 sky130_fd_sc_hd__nor2_4 _15587_ (.A(\CPU_Xreg_value_a4[26][6] ),
    .B(_09134_),
    .Y(_09225_));
 sky130_fd_sc_hd__a211o_4 _15588_ (.A1(_09224_),
    .A2(_09137_),
    .B1(_09215_),
    .C1(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__inv_2 _15589_ (.A(_09226_),
    .Y(_00180_));
 sky130_fd_sc_hd__buf_2 _15590_ (.A(_06837_),
    .X(_09227_));
 sky130_fd_sc_hd__nor2_4 _15591_ (.A(\CPU_Xreg_value_a4[26][5] ),
    .B(_09134_),
    .Y(_09228_));
 sky130_fd_sc_hd__a211o_4 _15592_ (.A1(_09227_),
    .A2(_09137_),
    .B1(_09215_),
    .C1(_09228_),
    .X(_09229_));
 sky130_fd_sc_hd__inv_2 _15593_ (.A(_09229_),
    .Y(_00179_));
 sky130_fd_sc_hd__buf_2 _15594_ (.A(_09134_),
    .X(_09230_));
 sky130_fd_sc_hd__inv_2 _15595_ (.A(\CPU_Xreg_value_a4[26][4] ),
    .Y(_09231_));
 sky130_fd_sc_hd__nor2_4 _15596_ (.A(_09231_),
    .B(_09230_),
    .Y(_09232_));
 sky130_fd_sc_hd__a211o_4 _15597_ (.A1(_08878_),
    .A2(_09230_),
    .B1(_09039_),
    .C1(_09232_),
    .X(_00178_));
 sky130_fd_sc_hd__buf_2 _15598_ (.A(_06102_),
    .X(_09233_));
 sky130_fd_sc_hd__inv_2 _15599_ (.A(\CPU_Xreg_value_a4[26][3] ),
    .Y(_09234_));
 sky130_fd_sc_hd__nor2_4 _15600_ (.A(_09234_),
    .B(_09230_),
    .Y(_09235_));
 sky130_fd_sc_hd__a211o_4 _15601_ (.A1(_08174_),
    .A2(_09230_),
    .B1(_09233_),
    .C1(_09235_),
    .X(_00177_));
 sky130_fd_sc_hd__nor2_4 _15602_ (.A(\CPU_Xreg_value_a4[26][2] ),
    .B(_09134_),
    .Y(_09236_));
 sky130_fd_sc_hd__a211o_4 _15603_ (.A1(_06860_),
    .A2(_09137_),
    .B1(_09215_),
    .C1(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__inv_2 _15604_ (.A(_09237_),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_2 _15605_ (.A(\CPU_Xreg_value_a4[26][1] ),
    .Y(_09238_));
 sky130_fd_sc_hd__nor2_4 _15606_ (.A(_09238_),
    .B(_09230_),
    .Y(_09239_));
 sky130_fd_sc_hd__a211o_4 _15607_ (.A1(_07096_),
    .A2(_09230_),
    .B1(_09233_),
    .C1(_09239_),
    .X(_00175_));
 sky130_fd_sc_hd__buf_2 _15608_ (.A(_09214_),
    .X(_09240_));
 sky130_fd_sc_hd__nor2_4 _15609_ (.A(\CPU_Xreg_value_a4[26][0] ),
    .B(_09134_),
    .Y(_09241_));
 sky130_fd_sc_hd__a211o_4 _15610_ (.A1(_07100_),
    .A2(_09137_),
    .B1(_09240_),
    .C1(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__inv_2 _15611_ (.A(_09242_),
    .Y(_00174_));
 sky130_fd_sc_hd__nor2_4 _15612_ (.A(_07821_),
    .B(_08362_),
    .Y(_09243_));
 sky130_fd_sc_hd__buf_2 _15613_ (.A(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__buf_2 _15614_ (.A(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__buf_2 _15615_ (.A(_09244_),
    .X(_09246_));
 sky130_fd_sc_hd__nor2_4 _15616_ (.A(\CPU_Xreg_value_a4[27][31] ),
    .B(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__a211o_4 _15617_ (.A1(_09132_),
    .A2(_09245_),
    .B1(_09240_),
    .C1(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__inv_2 _15618_ (.A(_09248_),
    .Y(_00173_));
 sky130_fd_sc_hd__nor2_4 _15619_ (.A(\CPU_Xreg_value_a4[27][30] ),
    .B(_09246_),
    .Y(_09249_));
 sky130_fd_sc_hd__a211o_4 _15620_ (.A1(_09140_),
    .A2(_09245_),
    .B1(_09240_),
    .C1(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__inv_2 _15621_ (.A(_09250_),
    .Y(_00172_));
 sky130_fd_sc_hd__nor2_4 _15622_ (.A(\CPU_Xreg_value_a4[27][29] ),
    .B(_09246_),
    .Y(_09251_));
 sky130_fd_sc_hd__a211o_4 _15623_ (.A1(_09144_),
    .A2(_09245_),
    .B1(_09240_),
    .C1(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__inv_2 _15624_ (.A(_09252_),
    .Y(_00171_));
 sky130_fd_sc_hd__nor2_4 _15625_ (.A(\CPU_Xreg_value_a4[27][28] ),
    .B(_09246_),
    .Y(_09253_));
 sky130_fd_sc_hd__a211o_4 _15626_ (.A1(_09147_),
    .A2(_09245_),
    .B1(_09240_),
    .C1(_09253_),
    .X(_09254_));
 sky130_fd_sc_hd__inv_2 _15627_ (.A(_09254_),
    .Y(_00170_));
 sky130_fd_sc_hd__buf_2 _15628_ (.A(_09243_),
    .X(_09255_));
 sky130_fd_sc_hd__buf_2 _15629_ (.A(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_4 _15630_ (.A(\CPU_Xreg_value_a4[27][27] ),
    .B(_09246_),
    .Y(_09257_));
 sky130_fd_sc_hd__a211o_4 _15631_ (.A1(_09150_),
    .A2(_09256_),
    .B1(_09240_),
    .C1(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__inv_2 _15632_ (.A(_09258_),
    .Y(_00169_));
 sky130_fd_sc_hd__buf_2 _15633_ (.A(_09214_),
    .X(_09259_));
 sky130_fd_sc_hd__nor2_4 _15634_ (.A(\CPU_Xreg_value_a4[27][26] ),
    .B(_09246_),
    .Y(_09260_));
 sky130_fd_sc_hd__a211o_4 _15635_ (.A1(_09154_),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__inv_2 _15636_ (.A(_09261_),
    .Y(_00168_));
 sky130_fd_sc_hd__buf_2 _15637_ (.A(_09244_),
    .X(_09262_));
 sky130_fd_sc_hd__nor2_4 _15638_ (.A(\CPU_Xreg_value_a4[27][25] ),
    .B(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__a211o_4 _15639_ (.A1(_09157_),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09263_),
    .X(_09264_));
 sky130_fd_sc_hd__inv_2 _15640_ (.A(_09264_),
    .Y(_00167_));
 sky130_fd_sc_hd__nor2_4 _15641_ (.A(\CPU_Xreg_value_a4[27][24] ),
    .B(_09262_),
    .Y(_09265_));
 sky130_fd_sc_hd__a211o_4 _15642_ (.A1(_09161_),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09265_),
    .X(_09266_));
 sky130_fd_sc_hd__inv_2 _15643_ (.A(_09266_),
    .Y(_00166_));
 sky130_fd_sc_hd__nor2_4 _15644_ (.A(\CPU_Xreg_value_a4[27][23] ),
    .B(_09262_),
    .Y(_09267_));
 sky130_fd_sc_hd__a211o_4 _15645_ (.A1(_09165_),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09267_),
    .X(_09268_));
 sky130_fd_sc_hd__inv_2 _15646_ (.A(_09268_),
    .Y(_00165_));
 sky130_fd_sc_hd__nor2_4 _15647_ (.A(\CPU_Xreg_value_a4[27][22] ),
    .B(_09262_),
    .Y(_09269_));
 sky130_fd_sc_hd__a211o_4 _15648_ (.A1(_09168_),
    .A2(_09256_),
    .B1(_09259_),
    .C1(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__inv_2 _15649_ (.A(_09270_),
    .Y(_00164_));
 sky130_fd_sc_hd__buf_2 _15650_ (.A(_09244_),
    .X(_09271_));
 sky130_fd_sc_hd__nor2_4 _15651_ (.A(\CPU_Xreg_value_a4[27][21] ),
    .B(_09262_),
    .Y(_09272_));
 sky130_fd_sc_hd__a211o_4 _15652_ (.A1(_09171_),
    .A2(_09271_),
    .B1(_09259_),
    .C1(_09272_),
    .X(_09273_));
 sky130_fd_sc_hd__inv_2 _15653_ (.A(_09273_),
    .Y(_00163_));
 sky130_fd_sc_hd__buf_2 _15654_ (.A(_09214_),
    .X(_09274_));
 sky130_fd_sc_hd__nor2_4 _15655_ (.A(\CPU_Xreg_value_a4[27][20] ),
    .B(_09262_),
    .Y(_09275_));
 sky130_fd_sc_hd__a211o_4 _15656_ (.A1(_09175_),
    .A2(_09271_),
    .B1(_09274_),
    .C1(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__inv_2 _15657_ (.A(_09276_),
    .Y(_00162_));
 sky130_fd_sc_hd__buf_2 _15658_ (.A(_09243_),
    .X(_09277_));
 sky130_fd_sc_hd__nor2_4 _15659_ (.A(\CPU_Xreg_value_a4[27][19] ),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__a211o_4 _15660_ (.A1(_09178_),
    .A2(_09271_),
    .B1(_09274_),
    .C1(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__inv_2 _15661_ (.A(_09279_),
    .Y(_00161_));
 sky130_fd_sc_hd__nor2_4 _15662_ (.A(\CPU_Xreg_value_a4[27][18] ),
    .B(_09277_),
    .Y(_09280_));
 sky130_fd_sc_hd__a211o_4 _15663_ (.A1(_09182_),
    .A2(_09271_),
    .B1(_09274_),
    .C1(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__inv_2 _15664_ (.A(_09281_),
    .Y(_00160_));
 sky130_fd_sc_hd__nor2_4 _15665_ (.A(\CPU_Xreg_value_a4[27][17] ),
    .B(_09277_),
    .Y(_09282_));
 sky130_fd_sc_hd__a211o_4 _15666_ (.A1(_09186_),
    .A2(_09271_),
    .B1(_09274_),
    .C1(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__inv_2 _15667_ (.A(_09283_),
    .Y(_00159_));
 sky130_fd_sc_hd__nor2_4 _15668_ (.A(\CPU_Xreg_value_a4[27][16] ),
    .B(_09277_),
    .Y(_09284_));
 sky130_fd_sc_hd__a211o_4 _15669_ (.A1(_09189_),
    .A2(_09271_),
    .B1(_09274_),
    .C1(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__inv_2 _15670_ (.A(_09285_),
    .Y(_00158_));
 sky130_fd_sc_hd__buf_2 _15671_ (.A(_09244_),
    .X(_09286_));
 sky130_fd_sc_hd__nor2_4 _15672_ (.A(\CPU_Xreg_value_a4[27][15] ),
    .B(_09277_),
    .Y(_09287_));
 sky130_fd_sc_hd__a211o_4 _15673_ (.A1(_09192_),
    .A2(_09286_),
    .B1(_09274_),
    .C1(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__inv_2 _15674_ (.A(_09288_),
    .Y(_00157_));
 sky130_fd_sc_hd__buf_2 _15675_ (.A(_09214_),
    .X(_09289_));
 sky130_fd_sc_hd__nor2_4 _15676_ (.A(\CPU_Xreg_value_a4[27][14] ),
    .B(_09277_),
    .Y(_09290_));
 sky130_fd_sc_hd__a211o_4 _15677_ (.A1(_09196_),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__inv_2 _15678_ (.A(_09291_),
    .Y(_00156_));
 sky130_fd_sc_hd__buf_2 _15679_ (.A(_09243_),
    .X(_09292_));
 sky130_fd_sc_hd__nor2_4 _15680_ (.A(\CPU_Xreg_value_a4[27][13] ),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a211o_4 _15681_ (.A1(_09199_),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__inv_2 _15682_ (.A(_09294_),
    .Y(_00155_));
 sky130_fd_sc_hd__nor2_4 _15683_ (.A(\CPU_Xreg_value_a4[27][12] ),
    .B(_09292_),
    .Y(_09295_));
 sky130_fd_sc_hd__a211o_4 _15684_ (.A1(_09203_),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09295_),
    .X(_09296_));
 sky130_fd_sc_hd__inv_2 _15685_ (.A(_09296_),
    .Y(_00154_));
 sky130_fd_sc_hd__nor2_4 _15686_ (.A(\CPU_Xreg_value_a4[27][11] ),
    .B(_09292_),
    .Y(_09297_));
 sky130_fd_sc_hd__a211o_4 _15687_ (.A1(_09207_),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__inv_2 _15688_ (.A(_09298_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2_4 _15689_ (.A(\CPU_Xreg_value_a4[27][10] ),
    .B(_09292_),
    .Y(_09299_));
 sky130_fd_sc_hd__a211o_4 _15690_ (.A1(_09210_),
    .A2(_09286_),
    .B1(_09289_),
    .C1(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__inv_2 _15691_ (.A(_09300_),
    .Y(_00152_));
 sky130_fd_sc_hd__buf_2 _15692_ (.A(_09244_),
    .X(_09301_));
 sky130_fd_sc_hd__nor2_4 _15693_ (.A(\CPU_Xreg_value_a4[27][9] ),
    .B(_09292_),
    .Y(_09302_));
 sky130_fd_sc_hd__a211o_4 _15694_ (.A1(_09213_),
    .A2(_09301_),
    .B1(_09289_),
    .C1(_09302_),
    .X(_09303_));
 sky130_fd_sc_hd__inv_2 _15695_ (.A(_09303_),
    .Y(_00151_));
 sky130_fd_sc_hd__buf_2 _15696_ (.A(_09214_),
    .X(_09304_));
 sky130_fd_sc_hd__nor2_4 _15697_ (.A(\CPU_Xreg_value_a4[27][8] ),
    .B(_09292_),
    .Y(_09305_));
 sky130_fd_sc_hd__a211o_4 _15698_ (.A1(_09218_),
    .A2(_09301_),
    .B1(_09304_),
    .C1(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__inv_2 _15699_ (.A(_09306_),
    .Y(_00150_));
 sky130_fd_sc_hd__nor2_4 _15700_ (.A(\CPU_Xreg_value_a4[27][7] ),
    .B(_09255_),
    .Y(_09307_));
 sky130_fd_sc_hd__a211o_4 _15701_ (.A1(_09221_),
    .A2(_09301_),
    .B1(_09304_),
    .C1(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__inv_2 _15702_ (.A(_09308_),
    .Y(_00149_));
 sky130_fd_sc_hd__nor2_4 _15703_ (.A(\CPU_Xreg_value_a4[27][6] ),
    .B(_09255_),
    .Y(_09309_));
 sky130_fd_sc_hd__a211o_4 _15704_ (.A1(_09224_),
    .A2(_09301_),
    .B1(_09304_),
    .C1(_09309_),
    .X(_09310_));
 sky130_fd_sc_hd__inv_2 _15705_ (.A(_09310_),
    .Y(_00148_));
 sky130_fd_sc_hd__nor2_4 _15706_ (.A(\CPU_Xreg_value_a4[27][5] ),
    .B(_09255_),
    .Y(_09311_));
 sky130_fd_sc_hd__a211o_4 _15707_ (.A1(_09227_),
    .A2(_09301_),
    .B1(_09304_),
    .C1(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__inv_2 _15708_ (.A(_09312_),
    .Y(_00147_));
 sky130_fd_sc_hd__buf_2 _15709_ (.A(_09255_),
    .X(_09313_));
 sky130_fd_sc_hd__inv_2 _15710_ (.A(\CPU_Xreg_value_a4[27][4] ),
    .Y(_09314_));
 sky130_fd_sc_hd__nor2_4 _15711_ (.A(_09314_),
    .B(_09313_),
    .Y(_09315_));
 sky130_fd_sc_hd__a211o_4 _15712_ (.A1(_08878_),
    .A2(_09313_),
    .B1(_09233_),
    .C1(_09315_),
    .X(_00146_));
 sky130_fd_sc_hd__inv_2 _15713_ (.A(\CPU_Xreg_value_a4[27][3] ),
    .Y(_09316_));
 sky130_fd_sc_hd__nor2_4 _15714_ (.A(_09316_),
    .B(_09313_),
    .Y(_09317_));
 sky130_fd_sc_hd__a211o_4 _15715_ (.A1(_08174_),
    .A2(_09313_),
    .B1(_09233_),
    .C1(_09317_),
    .X(_00145_));
 sky130_fd_sc_hd__nor2_4 _15716_ (.A(\CPU_Xreg_value_a4[27][2] ),
    .B(_09255_),
    .Y(_09318_));
 sky130_fd_sc_hd__a211o_4 _15717_ (.A1(_06860_),
    .A2(_09301_),
    .B1(_09304_),
    .C1(_09318_),
    .X(_09319_));
 sky130_fd_sc_hd__inv_2 _15718_ (.A(_09319_),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _15719_ (.A(\CPU_Xreg_value_a4[27][1] ),
    .Y(_09320_));
 sky130_fd_sc_hd__nor2_4 _15720_ (.A(_09320_),
    .B(_09245_),
    .Y(_09321_));
 sky130_fd_sc_hd__a211o_4 _15721_ (.A1(_07096_),
    .A2(_09313_),
    .B1(_09233_),
    .C1(_09321_),
    .X(_00143_));
 sky130_fd_sc_hd__inv_2 _15722_ (.A(\CPU_Xreg_value_a4[27][0] ),
    .Y(_09322_));
 sky130_fd_sc_hd__nor2_4 _15723_ (.A(_09322_),
    .B(_09245_),
    .Y(_09323_));
 sky130_fd_sc_hd__a211o_4 _15724_ (.A1(_06981_),
    .A2(_09313_),
    .B1(_09233_),
    .C1(_09323_),
    .X(_00142_));
 sky130_fd_sc_hd__or2_4 _15725_ (.A(_07905_),
    .B(_08362_),
    .X(_09324_));
 sky130_fd_sc_hd__inv_2 _15726_ (.A(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__buf_2 _15727_ (.A(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__buf_2 _15728_ (.A(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__buf_2 _15729_ (.A(_09325_),
    .X(_09328_));
 sky130_fd_sc_hd__nor2_4 _15730_ (.A(\CPU_Xreg_value_a4[28][31] ),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__a211o_4 _15731_ (.A1(_09132_),
    .A2(_09327_),
    .B1(_09304_),
    .C1(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__inv_2 _15732_ (.A(_09330_),
    .Y(_00141_));
 sky130_fd_sc_hd__buf_2 _15733_ (.A(_06100_),
    .X(_09331_));
 sky130_fd_sc_hd__buf_2 _15734_ (.A(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__nor2_4 _15735_ (.A(\CPU_Xreg_value_a4[28][30] ),
    .B(_09328_),
    .Y(_09333_));
 sky130_fd_sc_hd__a211o_4 _15736_ (.A1(_09140_),
    .A2(_09327_),
    .B1(_09332_),
    .C1(_09333_),
    .X(_09334_));
 sky130_fd_sc_hd__inv_2 _15737_ (.A(_09334_),
    .Y(_00140_));
 sky130_fd_sc_hd__nor2_4 _15738_ (.A(\CPU_Xreg_value_a4[28][29] ),
    .B(_09328_),
    .Y(_09335_));
 sky130_fd_sc_hd__a211o_4 _15739_ (.A1(_09144_),
    .A2(_09327_),
    .B1(_09332_),
    .C1(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__inv_2 _15740_ (.A(_09336_),
    .Y(_00139_));
 sky130_fd_sc_hd__buf_2 _15741_ (.A(_09326_),
    .X(_09337_));
 sky130_fd_sc_hd__nor2_4 _15742_ (.A(\CPU_Xreg_value_a4[28][28] ),
    .B(_09328_),
    .Y(_09338_));
 sky130_fd_sc_hd__a211o_4 _15743_ (.A1(_09147_),
    .A2(_09337_),
    .B1(_09332_),
    .C1(_09338_),
    .X(_09339_));
 sky130_fd_sc_hd__inv_2 _15744_ (.A(_09339_),
    .Y(_00138_));
 sky130_fd_sc_hd__buf_2 _15745_ (.A(_09325_),
    .X(_09340_));
 sky130_fd_sc_hd__nor2_4 _15746_ (.A(\CPU_Xreg_value_a4[28][27] ),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__a211o_4 _15747_ (.A1(_09150_),
    .A2(_09337_),
    .B1(_09332_),
    .C1(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__inv_2 _15748_ (.A(_09342_),
    .Y(_00137_));
 sky130_fd_sc_hd__nor2_4 _15749_ (.A(\CPU_Xreg_value_a4[28][26] ),
    .B(_09340_),
    .Y(_09343_));
 sky130_fd_sc_hd__a211o_4 _15750_ (.A1(_09154_),
    .A2(_09337_),
    .B1(_09332_),
    .C1(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__inv_2 _15751_ (.A(_09344_),
    .Y(_00136_));
 sky130_fd_sc_hd__nor2_4 _15752_ (.A(\CPU_Xreg_value_a4[28][25] ),
    .B(_09340_),
    .Y(_09345_));
 sky130_fd_sc_hd__a211o_4 _15753_ (.A1(_09157_),
    .A2(_09337_),
    .B1(_09332_),
    .C1(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__inv_2 _15754_ (.A(_09346_),
    .Y(_00135_));
 sky130_fd_sc_hd__buf_2 _15755_ (.A(_09331_),
    .X(_09347_));
 sky130_fd_sc_hd__nor2_4 _15756_ (.A(\CPU_Xreg_value_a4[28][24] ),
    .B(_09340_),
    .Y(_09348_));
 sky130_fd_sc_hd__a211o_4 _15757_ (.A1(_09161_),
    .A2(_09337_),
    .B1(_09347_),
    .C1(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__inv_2 _15758_ (.A(_09349_),
    .Y(_00134_));
 sky130_fd_sc_hd__nor2_4 _15759_ (.A(\CPU_Xreg_value_a4[28][23] ),
    .B(_09340_),
    .Y(_09350_));
 sky130_fd_sc_hd__a211o_4 _15760_ (.A1(_09165_),
    .A2(_09337_),
    .B1(_09347_),
    .C1(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__inv_2 _15761_ (.A(_09351_),
    .Y(_00133_));
 sky130_fd_sc_hd__buf_2 _15762_ (.A(_09326_),
    .X(_09352_));
 sky130_fd_sc_hd__nor2_4 _15763_ (.A(\CPU_Xreg_value_a4[28][22] ),
    .B(_09340_),
    .Y(_09353_));
 sky130_fd_sc_hd__a211o_4 _15764_ (.A1(_09168_),
    .A2(_09352_),
    .B1(_09347_),
    .C1(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__inv_2 _15765_ (.A(_09354_),
    .Y(_00132_));
 sky130_fd_sc_hd__buf_2 _15766_ (.A(_09325_),
    .X(_09355_));
 sky130_fd_sc_hd__nor2_4 _15767_ (.A(\CPU_Xreg_value_a4[28][21] ),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__a211o_4 _15768_ (.A1(_09171_),
    .A2(_09352_),
    .B1(_09347_),
    .C1(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__inv_2 _15769_ (.A(_09357_),
    .Y(_00131_));
 sky130_fd_sc_hd__nor2_4 _15770_ (.A(\CPU_Xreg_value_a4[28][20] ),
    .B(_09355_),
    .Y(_09358_));
 sky130_fd_sc_hd__a211o_4 _15771_ (.A1(_09175_),
    .A2(_09352_),
    .B1(_09347_),
    .C1(_09358_),
    .X(_09359_));
 sky130_fd_sc_hd__inv_2 _15772_ (.A(_09359_),
    .Y(_00130_));
 sky130_fd_sc_hd__nor2_4 _15773_ (.A(\CPU_Xreg_value_a4[28][19] ),
    .B(_09355_),
    .Y(_09360_));
 sky130_fd_sc_hd__a211o_4 _15774_ (.A1(_09178_),
    .A2(_09352_),
    .B1(_09347_),
    .C1(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__inv_2 _15775_ (.A(_09361_),
    .Y(_00129_));
 sky130_fd_sc_hd__buf_2 _15776_ (.A(_09331_),
    .X(_09362_));
 sky130_fd_sc_hd__nor2_4 _15777_ (.A(\CPU_Xreg_value_a4[28][18] ),
    .B(_09355_),
    .Y(_09363_));
 sky130_fd_sc_hd__a211o_4 _15778_ (.A1(_09182_),
    .A2(_09352_),
    .B1(_09362_),
    .C1(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__inv_2 _15779_ (.A(_09364_),
    .Y(_00128_));
 sky130_fd_sc_hd__nor2_4 _15780_ (.A(\CPU_Xreg_value_a4[28][17] ),
    .B(_09355_),
    .Y(_09365_));
 sky130_fd_sc_hd__a211o_4 _15781_ (.A1(_09186_),
    .A2(_09352_),
    .B1(_09362_),
    .C1(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__inv_2 _15782_ (.A(_09366_),
    .Y(_00127_));
 sky130_fd_sc_hd__buf_2 _15783_ (.A(_09326_),
    .X(_09367_));
 sky130_fd_sc_hd__nor2_4 _15784_ (.A(\CPU_Xreg_value_a4[28][16] ),
    .B(_09355_),
    .Y(_09368_));
 sky130_fd_sc_hd__a211o_4 _15785_ (.A1(_09189_),
    .A2(_09367_),
    .B1(_09362_),
    .C1(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__inv_2 _15786_ (.A(_09369_),
    .Y(_00126_));
 sky130_fd_sc_hd__buf_2 _15787_ (.A(_09325_),
    .X(_09370_));
 sky130_fd_sc_hd__nor2_4 _15788_ (.A(\CPU_Xreg_value_a4[28][15] ),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__a211o_4 _15789_ (.A1(_09192_),
    .A2(_09367_),
    .B1(_09362_),
    .C1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__inv_2 _15790_ (.A(_09372_),
    .Y(_00125_));
 sky130_fd_sc_hd__nor2_4 _15791_ (.A(\CPU_Xreg_value_a4[28][14] ),
    .B(_09370_),
    .Y(_09373_));
 sky130_fd_sc_hd__a211o_4 _15792_ (.A1(_09196_),
    .A2(_09367_),
    .B1(_09362_),
    .C1(_09373_),
    .X(_09374_));
 sky130_fd_sc_hd__inv_2 _15793_ (.A(_09374_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor2_4 _15794_ (.A(\CPU_Xreg_value_a4[28][13] ),
    .B(_09370_),
    .Y(_09375_));
 sky130_fd_sc_hd__a211o_4 _15795_ (.A1(_09199_),
    .A2(_09367_),
    .B1(_09362_),
    .C1(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__inv_2 _15796_ (.A(_09376_),
    .Y(_00123_));
 sky130_fd_sc_hd__buf_2 _15797_ (.A(_09331_),
    .X(_09377_));
 sky130_fd_sc_hd__nor2_4 _15798_ (.A(\CPU_Xreg_value_a4[28][12] ),
    .B(_09370_),
    .Y(_09378_));
 sky130_fd_sc_hd__a211o_4 _15799_ (.A1(_09203_),
    .A2(_09367_),
    .B1(_09377_),
    .C1(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__inv_2 _15800_ (.A(_09379_),
    .Y(_00122_));
 sky130_fd_sc_hd__nor2_4 _15801_ (.A(\CPU_Xreg_value_a4[28][11] ),
    .B(_09370_),
    .Y(_09380_));
 sky130_fd_sc_hd__a211o_4 _15802_ (.A1(_09207_),
    .A2(_09367_),
    .B1(_09377_),
    .C1(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__inv_2 _15803_ (.A(_09381_),
    .Y(_00121_));
 sky130_fd_sc_hd__buf_2 _15804_ (.A(_09326_),
    .X(_09382_));
 sky130_fd_sc_hd__nor2_4 _15805_ (.A(\CPU_Xreg_value_a4[28][10] ),
    .B(_09370_),
    .Y(_09383_));
 sky130_fd_sc_hd__a211o_4 _15806_ (.A1(_09210_),
    .A2(_09382_),
    .B1(_09377_),
    .C1(_09383_),
    .X(_09384_));
 sky130_fd_sc_hd__inv_2 _15807_ (.A(_09384_),
    .Y(_00120_));
 sky130_fd_sc_hd__buf_2 _15808_ (.A(_09325_),
    .X(_09385_));
 sky130_fd_sc_hd__nor2_4 _15809_ (.A(\CPU_Xreg_value_a4[28][9] ),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__a211o_4 _15810_ (.A1(_09213_),
    .A2(_09382_),
    .B1(_09377_),
    .C1(_09386_),
    .X(_09387_));
 sky130_fd_sc_hd__inv_2 _15811_ (.A(_09387_),
    .Y(_00119_));
 sky130_fd_sc_hd__nor2_4 _15812_ (.A(\CPU_Xreg_value_a4[28][8] ),
    .B(_09385_),
    .Y(_09388_));
 sky130_fd_sc_hd__a211o_4 _15813_ (.A1(_09218_),
    .A2(_09382_),
    .B1(_09377_),
    .C1(_09388_),
    .X(_09389_));
 sky130_fd_sc_hd__inv_2 _15814_ (.A(_09389_),
    .Y(_00118_));
 sky130_fd_sc_hd__nor2_4 _15815_ (.A(\CPU_Xreg_value_a4[28][7] ),
    .B(_09385_),
    .Y(_09390_));
 sky130_fd_sc_hd__a211o_4 _15816_ (.A1(_09221_),
    .A2(_09382_),
    .B1(_09377_),
    .C1(_09390_),
    .X(_09391_));
 sky130_fd_sc_hd__inv_2 _15817_ (.A(_09391_),
    .Y(_00117_));
 sky130_fd_sc_hd__buf_2 _15818_ (.A(_09331_),
    .X(_09392_));
 sky130_fd_sc_hd__nor2_4 _15819_ (.A(\CPU_Xreg_value_a4[28][6] ),
    .B(_09385_),
    .Y(_09393_));
 sky130_fd_sc_hd__a211o_4 _15820_ (.A1(_09224_),
    .A2(_09382_),
    .B1(_09392_),
    .C1(_09393_),
    .X(_09394_));
 sky130_fd_sc_hd__inv_2 _15821_ (.A(_09394_),
    .Y(_00116_));
 sky130_fd_sc_hd__nor2_4 _15822_ (.A(\CPU_Xreg_value_a4[28][5] ),
    .B(_09385_),
    .Y(_09395_));
 sky130_fd_sc_hd__a211o_4 _15823_ (.A1(_09227_),
    .A2(_09382_),
    .B1(_09392_),
    .C1(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__inv_2 _15824_ (.A(_09396_),
    .Y(_00115_));
 sky130_fd_sc_hd__buf_2 _15825_ (.A(_06102_),
    .X(_09397_));
 sky130_fd_sc_hd__and2_4 _15826_ (.A(\CPU_Xreg_value_a4[28][4] ),
    .B(_09324_),
    .X(_09398_));
 sky130_fd_sc_hd__a211o_4 _15827_ (.A1(_08345_),
    .A2(_09327_),
    .B1(_09397_),
    .C1(_09398_),
    .X(_00114_));
 sky130_fd_sc_hd__and2_4 _15828_ (.A(\CPU_Xreg_value_a4[28][3] ),
    .B(_09324_),
    .X(_09399_));
 sky130_fd_sc_hd__a211o_4 _15829_ (.A1(_07641_),
    .A2(_09327_),
    .B1(_09397_),
    .C1(_09399_),
    .X(_00113_));
 sky130_fd_sc_hd__and2_4 _15830_ (.A(\CPU_Xreg_value_a4[28][2] ),
    .B(_09324_),
    .X(_09400_));
 sky130_fd_sc_hd__a211o_4 _15831_ (.A1(_07271_),
    .A2(_09327_),
    .B1(_09397_),
    .C1(_09400_),
    .X(_00112_));
 sky130_fd_sc_hd__nor2_4 _15832_ (.A(\CPU_Xreg_value_a4[28][1] ),
    .B(_09385_),
    .Y(_09401_));
 sky130_fd_sc_hd__a211o_4 _15833_ (.A1(_06868_),
    .A2(_09328_),
    .B1(_09392_),
    .C1(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__inv_2 _15834_ (.A(_09402_),
    .Y(_00111_));
 sky130_fd_sc_hd__nor2_4 _15835_ (.A(\CPU_Xreg_value_a4[28][0] ),
    .B(_09326_),
    .Y(_09403_));
 sky130_fd_sc_hd__a211o_4 _15836_ (.A1(_07100_),
    .A2(_09328_),
    .B1(_09392_),
    .C1(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__inv_2 _15837_ (.A(_09404_),
    .Y(_00110_));
 sky130_fd_sc_hd__or2_4 _15838_ (.A(_07989_),
    .B(_08361_),
    .X(_09405_));
 sky130_fd_sc_hd__inv_2 _15839_ (.A(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__buf_2 _15840_ (.A(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__buf_2 _15841_ (.A(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__buf_2 _15842_ (.A(_09407_),
    .X(_09409_));
 sky130_fd_sc_hd__nor2_4 _15843_ (.A(\CPU_Xreg_value_a4[29][31] ),
    .B(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__a211o_4 _15844_ (.A1(_09132_),
    .A2(_09408_),
    .B1(_09392_),
    .C1(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__inv_2 _15845_ (.A(_09411_),
    .Y(_00109_));
 sky130_fd_sc_hd__nor2_4 _15846_ (.A(\CPU_Xreg_value_a4[29][30] ),
    .B(_09409_),
    .Y(_09412_));
 sky130_fd_sc_hd__a211o_4 _15847_ (.A1(_09140_),
    .A2(_09408_),
    .B1(_09392_),
    .C1(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__inv_2 _15848_ (.A(_09413_),
    .Y(_00108_));
 sky130_fd_sc_hd__buf_2 _15849_ (.A(_09407_),
    .X(_09414_));
 sky130_fd_sc_hd__buf_2 _15850_ (.A(_09331_),
    .X(_09415_));
 sky130_fd_sc_hd__nor2_4 _15851_ (.A(\CPU_Xreg_value_a4[29][29] ),
    .B(_09409_),
    .Y(_09416_));
 sky130_fd_sc_hd__a211o_4 _15852_ (.A1(_09144_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__inv_2 _15853_ (.A(_09417_),
    .Y(_00107_));
 sky130_fd_sc_hd__nor2_4 _15854_ (.A(\CPU_Xreg_value_a4[29][28] ),
    .B(_09409_),
    .Y(_09418_));
 sky130_fd_sc_hd__a211o_4 _15855_ (.A1(_09147_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__inv_2 _15856_ (.A(_09419_),
    .Y(_00106_));
 sky130_fd_sc_hd__buf_2 _15857_ (.A(_09406_),
    .X(_09420_));
 sky130_fd_sc_hd__nor2_4 _15858_ (.A(\CPU_Xreg_value_a4[29][27] ),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__a211o_4 _15859_ (.A1(_09150_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__inv_2 _15860_ (.A(_09422_),
    .Y(_00105_));
 sky130_fd_sc_hd__nor2_4 _15861_ (.A(\CPU_Xreg_value_a4[29][26] ),
    .B(_09420_),
    .Y(_09423_));
 sky130_fd_sc_hd__a211o_4 _15862_ (.A1(_09154_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__inv_2 _15863_ (.A(_09424_),
    .Y(_00104_));
 sky130_fd_sc_hd__nor2_4 _15864_ (.A(\CPU_Xreg_value_a4[29][25] ),
    .B(_09420_),
    .Y(_09425_));
 sky130_fd_sc_hd__a211o_4 _15865_ (.A1(_09157_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__inv_2 _15866_ (.A(_09426_),
    .Y(_00103_));
 sky130_fd_sc_hd__nor2_4 _15867_ (.A(\CPU_Xreg_value_a4[29][24] ),
    .B(_09420_),
    .Y(_09427_));
 sky130_fd_sc_hd__a211o_4 _15868_ (.A1(_09161_),
    .A2(_09414_),
    .B1(_09415_),
    .C1(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__inv_2 _15869_ (.A(_09428_),
    .Y(_00102_));
 sky130_fd_sc_hd__buf_2 _15870_ (.A(_09407_),
    .X(_09429_));
 sky130_fd_sc_hd__buf_2 _15871_ (.A(_06100_),
    .X(_09430_));
 sky130_fd_sc_hd__buf_2 _15872_ (.A(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__nor2_4 _15873_ (.A(\CPU_Xreg_value_a4[29][23] ),
    .B(_09420_),
    .Y(_09432_));
 sky130_fd_sc_hd__a211o_4 _15874_ (.A1(_09165_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__inv_2 _15875_ (.A(_09433_),
    .Y(_00101_));
 sky130_fd_sc_hd__nor2_4 _15876_ (.A(\CPU_Xreg_value_a4[29][22] ),
    .B(_09420_),
    .Y(_09434_));
 sky130_fd_sc_hd__a211o_4 _15877_ (.A1(_09168_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__inv_2 _15878_ (.A(_09435_),
    .Y(_00100_));
 sky130_fd_sc_hd__buf_2 _15879_ (.A(_09406_),
    .X(_09436_));
 sky130_fd_sc_hd__nor2_4 _15880_ (.A(\CPU_Xreg_value_a4[29][21] ),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__a211o_4 _15881_ (.A1(_09171_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09437_),
    .X(_09438_));
 sky130_fd_sc_hd__inv_2 _15882_ (.A(_09438_),
    .Y(_00099_));
 sky130_fd_sc_hd__nor2_4 _15883_ (.A(\CPU_Xreg_value_a4[29][20] ),
    .B(_09436_),
    .Y(_09439_));
 sky130_fd_sc_hd__a211o_4 _15884_ (.A1(_09175_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09439_),
    .X(_09440_));
 sky130_fd_sc_hd__inv_2 _15885_ (.A(_09440_),
    .Y(_00098_));
 sky130_fd_sc_hd__nor2_4 _15886_ (.A(\CPU_Xreg_value_a4[29][19] ),
    .B(_09436_),
    .Y(_09441_));
 sky130_fd_sc_hd__a211o_4 _15887_ (.A1(_09178_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__inv_2 _15888_ (.A(_09442_),
    .Y(_00097_));
 sky130_fd_sc_hd__nor2_4 _15889_ (.A(\CPU_Xreg_value_a4[29][18] ),
    .B(_09436_),
    .Y(_09443_));
 sky130_fd_sc_hd__a211o_4 _15890_ (.A1(_09182_),
    .A2(_09429_),
    .B1(_09431_),
    .C1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__inv_2 _15891_ (.A(_09444_),
    .Y(_00096_));
 sky130_fd_sc_hd__buf_2 _15892_ (.A(_09407_),
    .X(_09445_));
 sky130_fd_sc_hd__buf_2 _15893_ (.A(_09430_),
    .X(_09446_));
 sky130_fd_sc_hd__nor2_4 _15894_ (.A(\CPU_Xreg_value_a4[29][17] ),
    .B(_09436_),
    .Y(_09447_));
 sky130_fd_sc_hd__a211o_4 _15895_ (.A1(_09186_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__inv_2 _15896_ (.A(_09448_),
    .Y(_00095_));
 sky130_fd_sc_hd__nor2_4 _15897_ (.A(\CPU_Xreg_value_a4[29][16] ),
    .B(_09436_),
    .Y(_09449_));
 sky130_fd_sc_hd__a211o_4 _15898_ (.A1(_09189_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__inv_2 _15899_ (.A(_09450_),
    .Y(_00094_));
 sky130_fd_sc_hd__buf_2 _15900_ (.A(_09406_),
    .X(_09451_));
 sky130_fd_sc_hd__nor2_4 _15901_ (.A(\CPU_Xreg_value_a4[29][15] ),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__a211o_4 _15902_ (.A1(_09192_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09452_),
    .X(_09453_));
 sky130_fd_sc_hd__inv_2 _15903_ (.A(_09453_),
    .Y(_00093_));
 sky130_fd_sc_hd__nor2_4 _15904_ (.A(\CPU_Xreg_value_a4[29][14] ),
    .B(_09451_),
    .Y(_09454_));
 sky130_fd_sc_hd__a211o_4 _15905_ (.A1(_09196_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__inv_2 _15906_ (.A(_09455_),
    .Y(_00092_));
 sky130_fd_sc_hd__nor2_4 _15907_ (.A(\CPU_Xreg_value_a4[29][13] ),
    .B(_09451_),
    .Y(_09456_));
 sky130_fd_sc_hd__a211o_4 _15908_ (.A1(_09199_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09456_),
    .X(_09457_));
 sky130_fd_sc_hd__inv_2 _15909_ (.A(_09457_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor2_4 _15910_ (.A(\CPU_Xreg_value_a4[29][12] ),
    .B(_09451_),
    .Y(_09458_));
 sky130_fd_sc_hd__a211o_4 _15911_ (.A1(_09203_),
    .A2(_09445_),
    .B1(_09446_),
    .C1(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__inv_2 _15912_ (.A(_09459_),
    .Y(_00090_));
 sky130_fd_sc_hd__buf_2 _15913_ (.A(_09407_),
    .X(_09460_));
 sky130_fd_sc_hd__buf_2 _15914_ (.A(_09430_),
    .X(_09461_));
 sky130_fd_sc_hd__nor2_4 _15915_ (.A(\CPU_Xreg_value_a4[29][11] ),
    .B(_09451_),
    .Y(_09462_));
 sky130_fd_sc_hd__a211o_4 _15916_ (.A1(_09207_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__inv_2 _15917_ (.A(_09463_),
    .Y(_00089_));
 sky130_fd_sc_hd__nor2_4 _15918_ (.A(\CPU_Xreg_value_a4[29][10] ),
    .B(_09451_),
    .Y(_09464_));
 sky130_fd_sc_hd__a211o_4 _15919_ (.A1(_09210_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__inv_2 _15920_ (.A(_09465_),
    .Y(_00088_));
 sky130_fd_sc_hd__buf_2 _15921_ (.A(_09406_),
    .X(_09466_));
 sky130_fd_sc_hd__nor2_4 _15922_ (.A(\CPU_Xreg_value_a4[29][9] ),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__a211o_4 _15923_ (.A1(_09213_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__inv_2 _15924_ (.A(_09468_),
    .Y(_00087_));
 sky130_fd_sc_hd__nor2_4 _15925_ (.A(\CPU_Xreg_value_a4[29][8] ),
    .B(_09466_),
    .Y(_09469_));
 sky130_fd_sc_hd__a211o_4 _15926_ (.A1(_09218_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__inv_2 _15927_ (.A(_09470_),
    .Y(_00086_));
 sky130_fd_sc_hd__nor2_4 _15928_ (.A(\CPU_Xreg_value_a4[29][7] ),
    .B(_09466_),
    .Y(_09471_));
 sky130_fd_sc_hd__a211o_4 _15929_ (.A1(_09221_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__inv_2 _15930_ (.A(_09472_),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2_4 _15931_ (.A(\CPU_Xreg_value_a4[29][6] ),
    .B(_09466_),
    .Y(_09473_));
 sky130_fd_sc_hd__a211o_4 _15932_ (.A1(_09224_),
    .A2(_09460_),
    .B1(_09461_),
    .C1(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__inv_2 _15933_ (.A(_09474_),
    .Y(_00084_));
 sky130_fd_sc_hd__buf_2 _15934_ (.A(_09430_),
    .X(_09475_));
 sky130_fd_sc_hd__nor2_4 _15935_ (.A(\CPU_Xreg_value_a4[29][5] ),
    .B(_09466_),
    .Y(_09476_));
 sky130_fd_sc_hd__a211o_4 _15936_ (.A1(_09227_),
    .A2(_09409_),
    .B1(_09475_),
    .C1(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__inv_2 _15937_ (.A(_09477_),
    .Y(_00083_));
 sky130_fd_sc_hd__and2_4 _15938_ (.A(\CPU_Xreg_value_a4[29][4] ),
    .B(_09405_),
    .X(_09478_));
 sky130_fd_sc_hd__a211o_4 _15939_ (.A1(_08345_),
    .A2(_09408_),
    .B1(_09397_),
    .C1(_09478_),
    .X(_00082_));
 sky130_fd_sc_hd__and2_4 _15940_ (.A(\CPU_Xreg_value_a4[29][3] ),
    .B(_09405_),
    .X(_09479_));
 sky130_fd_sc_hd__a211o_4 _15941_ (.A1(_07641_),
    .A2(_09408_),
    .B1(_09397_),
    .C1(_09479_),
    .X(_00081_));
 sky130_fd_sc_hd__and2_4 _15942_ (.A(\CPU_Xreg_value_a4[29][2] ),
    .B(_09405_),
    .X(_09480_));
 sky130_fd_sc_hd__a211o_4 _15943_ (.A1(_07271_),
    .A2(_09408_),
    .B1(_09397_),
    .C1(_09480_),
    .X(_00080_));
 sky130_fd_sc_hd__nor2_4 _15944_ (.A(\CPU_Xreg_value_a4[29][1] ),
    .B(_09466_),
    .Y(_09481_));
 sky130_fd_sc_hd__a211o_4 _15945_ (.A1(_06868_),
    .A2(_09409_),
    .B1(_09475_),
    .C1(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__inv_2 _15946_ (.A(_09482_),
    .Y(_00079_));
 sky130_fd_sc_hd__buf_2 _15947_ (.A(_06102_),
    .X(_09483_));
 sky130_fd_sc_hd__and2_4 _15948_ (.A(\CPU_Xreg_value_a4[29][0] ),
    .B(_09405_),
    .X(_09484_));
 sky130_fd_sc_hd__a211o_4 _15949_ (.A1(_06981_),
    .A2(_09408_),
    .B1(_09483_),
    .C1(_09484_),
    .X(_00078_));
 sky130_fd_sc_hd__or2_4 _15950_ (.A(_08073_),
    .B(_08361_),
    .X(_09485_));
 sky130_fd_sc_hd__inv_2 _15951_ (.A(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__buf_2 _15952_ (.A(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__buf_2 _15953_ (.A(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__buf_2 _15954_ (.A(_09487_),
    .X(_09489_));
 sky130_fd_sc_hd__nor2_4 _15955_ (.A(\CPU_Xreg_value_a4[30][31] ),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__a211o_4 _15956_ (.A1(_09132_),
    .A2(_09488_),
    .B1(_09475_),
    .C1(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__inv_2 _15957_ (.A(_09491_),
    .Y(_00077_));
 sky130_fd_sc_hd__nor2_4 _15958_ (.A(\CPU_Xreg_value_a4[30][30] ),
    .B(_09489_),
    .Y(_09492_));
 sky130_fd_sc_hd__a211o_4 _15959_ (.A1(_09140_),
    .A2(_09488_),
    .B1(_09475_),
    .C1(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__inv_2 _15960_ (.A(_09493_),
    .Y(_00076_));
 sky130_fd_sc_hd__buf_2 _15961_ (.A(_09487_),
    .X(_09494_));
 sky130_fd_sc_hd__nor2_4 _15962_ (.A(\CPU_Xreg_value_a4[30][29] ),
    .B(_09489_),
    .Y(_09495_));
 sky130_fd_sc_hd__a211o_4 _15963_ (.A1(_09144_),
    .A2(_09494_),
    .B1(_09475_),
    .C1(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__inv_2 _15964_ (.A(_09496_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor2_4 _15965_ (.A(\CPU_Xreg_value_a4[30][28] ),
    .B(_09489_),
    .Y(_09497_));
 sky130_fd_sc_hd__a211o_4 _15966_ (.A1(_09147_),
    .A2(_09494_),
    .B1(_09475_),
    .C1(_09497_),
    .X(_09498_));
 sky130_fd_sc_hd__inv_2 _15967_ (.A(_09498_),
    .Y(_00074_));
 sky130_fd_sc_hd__buf_2 _15968_ (.A(_09430_),
    .X(_09499_));
 sky130_fd_sc_hd__buf_2 _15969_ (.A(_09486_),
    .X(_09500_));
 sky130_fd_sc_hd__nor2_4 _15970_ (.A(\CPU_Xreg_value_a4[30][27] ),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__a211o_4 _15971_ (.A1(_09150_),
    .A2(_09494_),
    .B1(_09499_),
    .C1(_09501_),
    .X(_09502_));
 sky130_fd_sc_hd__inv_2 _15972_ (.A(_09502_),
    .Y(_00073_));
 sky130_fd_sc_hd__nor2_4 _15973_ (.A(\CPU_Xreg_value_a4[30][26] ),
    .B(_09500_),
    .Y(_09503_));
 sky130_fd_sc_hd__a211o_4 _15974_ (.A1(_09154_),
    .A2(_09494_),
    .B1(_09499_),
    .C1(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__inv_2 _15975_ (.A(_09504_),
    .Y(_00072_));
 sky130_fd_sc_hd__nor2_4 _15976_ (.A(\CPU_Xreg_value_a4[30][25] ),
    .B(_09500_),
    .Y(_09505_));
 sky130_fd_sc_hd__a211o_4 _15977_ (.A1(_09157_),
    .A2(_09494_),
    .B1(_09499_),
    .C1(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__inv_2 _15978_ (.A(_09506_),
    .Y(_00071_));
 sky130_fd_sc_hd__nor2_4 _15979_ (.A(\CPU_Xreg_value_a4[30][24] ),
    .B(_09500_),
    .Y(_09507_));
 sky130_fd_sc_hd__a211o_4 _15980_ (.A1(_09161_),
    .A2(_09494_),
    .B1(_09499_),
    .C1(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__inv_2 _15981_ (.A(_09508_),
    .Y(_00070_));
 sky130_fd_sc_hd__buf_2 _15982_ (.A(_09487_),
    .X(_09509_));
 sky130_fd_sc_hd__nor2_4 _15983_ (.A(\CPU_Xreg_value_a4[30][23] ),
    .B(_09500_),
    .Y(_09510_));
 sky130_fd_sc_hd__a211o_4 _15984_ (.A1(_09165_),
    .A2(_09509_),
    .B1(_09499_),
    .C1(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__inv_2 _15985_ (.A(_09511_),
    .Y(_00069_));
 sky130_fd_sc_hd__nor2_4 _15986_ (.A(\CPU_Xreg_value_a4[30][22] ),
    .B(_09500_),
    .Y(_09512_));
 sky130_fd_sc_hd__a211o_4 _15987_ (.A1(_09168_),
    .A2(_09509_),
    .B1(_09499_),
    .C1(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__inv_2 _15988_ (.A(_09513_),
    .Y(_00068_));
 sky130_fd_sc_hd__buf_2 _15989_ (.A(_09430_),
    .X(_09514_));
 sky130_fd_sc_hd__buf_2 _15990_ (.A(_09486_),
    .X(_09515_));
 sky130_fd_sc_hd__nor2_4 _15991_ (.A(\CPU_Xreg_value_a4[30][21] ),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__a211o_4 _15992_ (.A1(_09171_),
    .A2(_09509_),
    .B1(_09514_),
    .C1(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__inv_2 _15993_ (.A(_09517_),
    .Y(_00067_));
 sky130_fd_sc_hd__nor2_4 _15994_ (.A(\CPU_Xreg_value_a4[30][20] ),
    .B(_09515_),
    .Y(_09518_));
 sky130_fd_sc_hd__a211o_4 _15995_ (.A1(_09175_),
    .A2(_09509_),
    .B1(_09514_),
    .C1(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__inv_2 _15996_ (.A(_09519_),
    .Y(_00066_));
 sky130_fd_sc_hd__nor2_4 _15997_ (.A(\CPU_Xreg_value_a4[30][19] ),
    .B(_09515_),
    .Y(_09520_));
 sky130_fd_sc_hd__a211o_4 _15998_ (.A1(_09178_),
    .A2(_09509_),
    .B1(_09514_),
    .C1(_09520_),
    .X(_09521_));
 sky130_fd_sc_hd__inv_2 _15999_ (.A(_09521_),
    .Y(_00065_));
 sky130_fd_sc_hd__nor2_4 _16000_ (.A(\CPU_Xreg_value_a4[30][18] ),
    .B(_09515_),
    .Y(_09522_));
 sky130_fd_sc_hd__a211o_4 _16001_ (.A1(_09182_),
    .A2(_09509_),
    .B1(_09514_),
    .C1(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__inv_2 _16002_ (.A(_09523_),
    .Y(_00064_));
 sky130_fd_sc_hd__buf_2 _16003_ (.A(_09487_),
    .X(_09524_));
 sky130_fd_sc_hd__nor2_4 _16004_ (.A(\CPU_Xreg_value_a4[30][17] ),
    .B(_09515_),
    .Y(_09525_));
 sky130_fd_sc_hd__a211o_4 _16005_ (.A1(_09186_),
    .A2(_09524_),
    .B1(_09514_),
    .C1(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__inv_2 _16006_ (.A(_09526_),
    .Y(_00063_));
 sky130_fd_sc_hd__nor2_4 _16007_ (.A(\CPU_Xreg_value_a4[30][16] ),
    .B(_09515_),
    .Y(_09527_));
 sky130_fd_sc_hd__a211o_4 _16008_ (.A1(_09189_),
    .A2(_09524_),
    .B1(_09514_),
    .C1(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__inv_2 _16009_ (.A(_09528_),
    .Y(_00062_));
 sky130_fd_sc_hd__buf_2 _16010_ (.A(_06100_),
    .X(_09529_));
 sky130_fd_sc_hd__buf_2 _16011_ (.A(_09529_),
    .X(_09530_));
 sky130_fd_sc_hd__buf_2 _16012_ (.A(_09486_),
    .X(_09531_));
 sky130_fd_sc_hd__nor2_4 _16013_ (.A(\CPU_Xreg_value_a4[30][15] ),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__a211o_4 _16014_ (.A1(_09192_),
    .A2(_09524_),
    .B1(_09530_),
    .C1(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__inv_2 _16015_ (.A(_09533_),
    .Y(_00061_));
 sky130_fd_sc_hd__nor2_4 _16016_ (.A(\CPU_Xreg_value_a4[30][14] ),
    .B(_09531_),
    .Y(_09534_));
 sky130_fd_sc_hd__a211o_4 _16017_ (.A1(_09196_),
    .A2(_09524_),
    .B1(_09530_),
    .C1(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__inv_2 _16018_ (.A(_09535_),
    .Y(_00060_));
 sky130_fd_sc_hd__nor2_4 _16019_ (.A(\CPU_Xreg_value_a4[30][13] ),
    .B(_09531_),
    .Y(_09536_));
 sky130_fd_sc_hd__a211o_4 _16020_ (.A1(_09199_),
    .A2(_09524_),
    .B1(_09530_),
    .C1(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__inv_2 _16021_ (.A(_09537_),
    .Y(_00059_));
 sky130_fd_sc_hd__nor2_4 _16022_ (.A(\CPU_Xreg_value_a4[30][12] ),
    .B(_09531_),
    .Y(_09538_));
 sky130_fd_sc_hd__a211o_4 _16023_ (.A1(_09203_),
    .A2(_09524_),
    .B1(_09530_),
    .C1(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__inv_2 _16024_ (.A(_09539_),
    .Y(_00058_));
 sky130_fd_sc_hd__buf_2 _16025_ (.A(_09487_),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_4 _16026_ (.A(\CPU_Xreg_value_a4[30][11] ),
    .B(_09531_),
    .Y(_09541_));
 sky130_fd_sc_hd__a211o_4 _16027_ (.A1(_09207_),
    .A2(_09540_),
    .B1(_09530_),
    .C1(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__inv_2 _16028_ (.A(_09542_),
    .Y(_00057_));
 sky130_fd_sc_hd__nor2_4 _16029_ (.A(\CPU_Xreg_value_a4[30][10] ),
    .B(_09531_),
    .Y(_09543_));
 sky130_fd_sc_hd__a211o_4 _16030_ (.A1(_09210_),
    .A2(_09540_),
    .B1(_09530_),
    .C1(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__inv_2 _16031_ (.A(_09544_),
    .Y(_00056_));
 sky130_fd_sc_hd__buf_2 _16032_ (.A(_09529_),
    .X(_09545_));
 sky130_fd_sc_hd__buf_2 _16033_ (.A(_09486_),
    .X(_09546_));
 sky130_fd_sc_hd__nor2_4 _16034_ (.A(\CPU_Xreg_value_a4[30][9] ),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__a211o_4 _16035_ (.A1(_09213_),
    .A2(_09540_),
    .B1(_09545_),
    .C1(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__inv_2 _16036_ (.A(_09548_),
    .Y(_00055_));
 sky130_fd_sc_hd__nor2_4 _16037_ (.A(\CPU_Xreg_value_a4[30][8] ),
    .B(_09546_),
    .Y(_09549_));
 sky130_fd_sc_hd__a211o_4 _16038_ (.A1(_09218_),
    .A2(_09540_),
    .B1(_09545_),
    .C1(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__inv_2 _16039_ (.A(_09550_),
    .Y(_00054_));
 sky130_fd_sc_hd__nor2_4 _16040_ (.A(\CPU_Xreg_value_a4[30][7] ),
    .B(_09546_),
    .Y(_09551_));
 sky130_fd_sc_hd__a211o_4 _16041_ (.A1(_09221_),
    .A2(_09540_),
    .B1(_09545_),
    .C1(_09551_),
    .X(_09552_));
 sky130_fd_sc_hd__inv_2 _16042_ (.A(_09552_),
    .Y(_00053_));
 sky130_fd_sc_hd__nor2_4 _16043_ (.A(\CPU_Xreg_value_a4[30][6] ),
    .B(_09546_),
    .Y(_09553_));
 sky130_fd_sc_hd__a211o_4 _16044_ (.A1(_09224_),
    .A2(_09540_),
    .B1(_09545_),
    .C1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__inv_2 _16045_ (.A(_09554_),
    .Y(_00052_));
 sky130_fd_sc_hd__nor2_4 _16046_ (.A(\CPU_Xreg_value_a4[30][5] ),
    .B(_09546_),
    .Y(_09555_));
 sky130_fd_sc_hd__a211o_4 _16047_ (.A1(_09227_),
    .A2(_09489_),
    .B1(_09545_),
    .C1(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__inv_2 _16048_ (.A(_09556_),
    .Y(_00051_));
 sky130_fd_sc_hd__and2_4 _16049_ (.A(\CPU_Xreg_value_a4[30][4] ),
    .B(_09485_),
    .X(_09557_));
 sky130_fd_sc_hd__a211o_4 _16050_ (.A1(_08345_),
    .A2(_09488_),
    .B1(_09483_),
    .C1(_09557_),
    .X(_00050_));
 sky130_fd_sc_hd__and2_4 _16051_ (.A(\CPU_Xreg_value_a4[30][3] ),
    .B(_09485_),
    .X(_09558_));
 sky130_fd_sc_hd__a211o_4 _16052_ (.A1(_07641_),
    .A2(_09488_),
    .B1(_09483_),
    .C1(_09558_),
    .X(_00049_));
 sky130_fd_sc_hd__and2_4 _16053_ (.A(\CPU_Xreg_value_a4[30][2] ),
    .B(_09485_),
    .X(_09559_));
 sky130_fd_sc_hd__a211o_4 _16054_ (.A1(_07271_),
    .A2(_09488_),
    .B1(_09483_),
    .C1(_09559_),
    .X(_00048_));
 sky130_fd_sc_hd__and2_4 _16055_ (.A(\CPU_Xreg_value_a4[30][1] ),
    .B(_09485_),
    .X(_09560_));
 sky130_fd_sc_hd__a211o_4 _16056_ (.A1(_07096_),
    .A2(_09488_),
    .B1(_09483_),
    .C1(_09560_),
    .X(_00047_));
 sky130_fd_sc_hd__nor2_4 _16057_ (.A(\CPU_Xreg_value_a4[30][0] ),
    .B(_09546_),
    .Y(_09561_));
 sky130_fd_sc_hd__a211o_4 _16058_ (.A1(_07100_),
    .A2(_09489_),
    .B1(_09545_),
    .C1(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__inv_2 _16059_ (.A(_09562_),
    .Y(_00046_));
 sky130_fd_sc_hd__or2_4 _16060_ (.A(_08187_),
    .B(_08361_),
    .X(_09563_));
 sky130_fd_sc_hd__inv_2 _16061_ (.A(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__buf_2 _16062_ (.A(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__buf_2 _16063_ (.A(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__buf_2 _16064_ (.A(_09529_),
    .X(_09567_));
 sky130_fd_sc_hd__buf_2 _16065_ (.A(_09564_),
    .X(_09568_));
 sky130_fd_sc_hd__buf_2 _16066_ (.A(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__nor2_4 _16067_ (.A(\CPU_Xreg_value_a4[31][31] ),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__a211o_4 _16068_ (.A1(_09132_),
    .A2(_09566_),
    .B1(_09567_),
    .C1(_09570_),
    .X(_09571_));
 sky130_fd_sc_hd__inv_2 _16069_ (.A(_09571_),
    .Y(_00045_));
 sky130_fd_sc_hd__buf_2 _16070_ (.A(_09568_),
    .X(_09572_));
 sky130_fd_sc_hd__nor2_4 _16071_ (.A(\CPU_Xreg_value_a4[31][30] ),
    .B(_09569_),
    .Y(_09573_));
 sky130_fd_sc_hd__a211o_4 _16072_ (.A1(_09140_),
    .A2(_09572_),
    .B1(_09567_),
    .C1(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__inv_2 _16073_ (.A(_09574_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_4 _16074_ (.A(\CPU_Xreg_value_a4[31][29] ),
    .B(_09569_),
    .Y(_09575_));
 sky130_fd_sc_hd__a211o_4 _16075_ (.A1(_09144_),
    .A2(_09572_),
    .B1(_09567_),
    .C1(_09575_),
    .X(_09576_));
 sky130_fd_sc_hd__inv_2 _16076_ (.A(_09576_),
    .Y(_00043_));
 sky130_fd_sc_hd__nor2_4 _16077_ (.A(\CPU_Xreg_value_a4[31][28] ),
    .B(_09569_),
    .Y(_09577_));
 sky130_fd_sc_hd__a211o_4 _16078_ (.A1(_09147_),
    .A2(_09572_),
    .B1(_09567_),
    .C1(_09577_),
    .X(_09578_));
 sky130_fd_sc_hd__inv_2 _16079_ (.A(_09578_),
    .Y(_00042_));
 sky130_fd_sc_hd__buf_2 _16080_ (.A(_09568_),
    .X(_09579_));
 sky130_fd_sc_hd__nor2_4 _16081_ (.A(\CPU_Xreg_value_a4[31][27] ),
    .B(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__a211o_4 _16082_ (.A1(_09150_),
    .A2(_09572_),
    .B1(_09567_),
    .C1(_09580_),
    .X(_09581_));
 sky130_fd_sc_hd__inv_2 _16083_ (.A(_09581_),
    .Y(_00041_));
 sky130_fd_sc_hd__nor2_4 _16084_ (.A(\CPU_Xreg_value_a4[31][26] ),
    .B(_09579_),
    .Y(_09582_));
 sky130_fd_sc_hd__a211o_4 _16085_ (.A1(_09154_),
    .A2(_09572_),
    .B1(_09567_),
    .C1(_09582_),
    .X(_09583_));
 sky130_fd_sc_hd__inv_2 _16086_ (.A(_09583_),
    .Y(_00040_));
 sky130_fd_sc_hd__buf_2 _16087_ (.A(_09529_),
    .X(_09584_));
 sky130_fd_sc_hd__nor2_4 _16088_ (.A(\CPU_Xreg_value_a4[31][25] ),
    .B(_09579_),
    .Y(_09585_));
 sky130_fd_sc_hd__a211o_4 _16089_ (.A1(_09157_),
    .A2(_09572_),
    .B1(_09584_),
    .C1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__inv_2 _16090_ (.A(_09586_),
    .Y(_00039_));
 sky130_fd_sc_hd__buf_2 _16091_ (.A(_09568_),
    .X(_09587_));
 sky130_fd_sc_hd__nor2_4 _16092_ (.A(\CPU_Xreg_value_a4[31][24] ),
    .B(_09579_),
    .Y(_09588_));
 sky130_fd_sc_hd__a211o_4 _16093_ (.A1(_09161_),
    .A2(_09587_),
    .B1(_09584_),
    .C1(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__inv_2 _16094_ (.A(_09589_),
    .Y(_00038_));
 sky130_fd_sc_hd__nor2_4 _16095_ (.A(\CPU_Xreg_value_a4[31][23] ),
    .B(_09579_),
    .Y(_09590_));
 sky130_fd_sc_hd__a211o_4 _16096_ (.A1(_09165_),
    .A2(_09587_),
    .B1(_09584_),
    .C1(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__inv_2 _16097_ (.A(_09591_),
    .Y(_00037_));
 sky130_fd_sc_hd__nor2_4 _16098_ (.A(\CPU_Xreg_value_a4[31][22] ),
    .B(_09579_),
    .Y(_09592_));
 sky130_fd_sc_hd__a211o_4 _16099_ (.A1(_09168_),
    .A2(_09587_),
    .B1(_09584_),
    .C1(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__inv_2 _16100_ (.A(_09593_),
    .Y(_00036_));
 sky130_fd_sc_hd__buf_2 _16101_ (.A(_09564_),
    .X(_09594_));
 sky130_fd_sc_hd__nor2_4 _16102_ (.A(\CPU_Xreg_value_a4[31][21] ),
    .B(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__a211o_4 _16103_ (.A1(_09171_),
    .A2(_09587_),
    .B1(_09584_),
    .C1(_09595_),
    .X(_09596_));
 sky130_fd_sc_hd__inv_2 _16104_ (.A(_09596_),
    .Y(_00035_));
 sky130_fd_sc_hd__nor2_4 _16105_ (.A(\CPU_Xreg_value_a4[31][20] ),
    .B(_09594_),
    .Y(_09597_));
 sky130_fd_sc_hd__a211o_4 _16106_ (.A1(_09175_),
    .A2(_09587_),
    .B1(_09584_),
    .C1(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__inv_2 _16107_ (.A(_09598_),
    .Y(_00034_));
 sky130_fd_sc_hd__buf_2 _16108_ (.A(_09529_),
    .X(_09599_));
 sky130_fd_sc_hd__nor2_4 _16109_ (.A(\CPU_Xreg_value_a4[31][19] ),
    .B(_09594_),
    .Y(_09600_));
 sky130_fd_sc_hd__a211o_4 _16110_ (.A1(_09178_),
    .A2(_09587_),
    .B1(_09599_),
    .C1(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__inv_2 _16111_ (.A(_09601_),
    .Y(_00033_));
 sky130_fd_sc_hd__buf_2 _16112_ (.A(_09568_),
    .X(_09602_));
 sky130_fd_sc_hd__nor2_4 _16113_ (.A(\CPU_Xreg_value_a4[31][18] ),
    .B(_09594_),
    .Y(_09603_));
 sky130_fd_sc_hd__a211o_4 _16114_ (.A1(_09182_),
    .A2(_09602_),
    .B1(_09599_),
    .C1(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__inv_2 _16115_ (.A(_09604_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_4 _16116_ (.A(\CPU_Xreg_value_a4[31][17] ),
    .B(_09594_),
    .Y(_09605_));
 sky130_fd_sc_hd__a211o_4 _16117_ (.A1(_09186_),
    .A2(_09602_),
    .B1(_09599_),
    .C1(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__inv_2 _16118_ (.A(_09606_),
    .Y(_00031_));
 sky130_fd_sc_hd__nor2_4 _16119_ (.A(\CPU_Xreg_value_a4[31][16] ),
    .B(_09594_),
    .Y(_09607_));
 sky130_fd_sc_hd__a211o_4 _16120_ (.A1(_09189_),
    .A2(_09602_),
    .B1(_09599_),
    .C1(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__inv_2 _16121_ (.A(_09608_),
    .Y(_00030_));
 sky130_fd_sc_hd__buf_2 _16122_ (.A(_09564_),
    .X(_09609_));
 sky130_fd_sc_hd__nor2_4 _16123_ (.A(\CPU_Xreg_value_a4[31][15] ),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__a211o_4 _16124_ (.A1(_09192_),
    .A2(_09602_),
    .B1(_09599_),
    .C1(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__inv_2 _16125_ (.A(_09611_),
    .Y(_00029_));
 sky130_fd_sc_hd__nor2_4 _16126_ (.A(\CPU_Xreg_value_a4[31][14] ),
    .B(_09609_),
    .Y(_09612_));
 sky130_fd_sc_hd__a211o_4 _16127_ (.A1(_09196_),
    .A2(_09602_),
    .B1(_09599_),
    .C1(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__inv_2 _16128_ (.A(_09613_),
    .Y(_00028_));
 sky130_fd_sc_hd__buf_2 _16129_ (.A(_09529_),
    .X(_09614_));
 sky130_fd_sc_hd__nor2_4 _16130_ (.A(\CPU_Xreg_value_a4[31][13] ),
    .B(_09609_),
    .Y(_09615_));
 sky130_fd_sc_hd__a211o_4 _16131_ (.A1(_09199_),
    .A2(_09602_),
    .B1(_09614_),
    .C1(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__inv_2 _16132_ (.A(_09616_),
    .Y(_00027_));
 sky130_fd_sc_hd__buf_2 _16133_ (.A(_09568_),
    .X(_09617_));
 sky130_fd_sc_hd__nor2_4 _16134_ (.A(\CPU_Xreg_value_a4[31][12] ),
    .B(_09609_),
    .Y(_09618_));
 sky130_fd_sc_hd__a211o_4 _16135_ (.A1(_09203_),
    .A2(_09617_),
    .B1(_09614_),
    .C1(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__inv_2 _16136_ (.A(_09619_),
    .Y(_00026_));
 sky130_fd_sc_hd__nor2_4 _16137_ (.A(\CPU_Xreg_value_a4[31][11] ),
    .B(_09609_),
    .Y(_09620_));
 sky130_fd_sc_hd__a211o_4 _16138_ (.A1(_09207_),
    .A2(_09617_),
    .B1(_09614_),
    .C1(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__inv_2 _16139_ (.A(_09621_),
    .Y(_00025_));
 sky130_fd_sc_hd__nor2_4 _16140_ (.A(\CPU_Xreg_value_a4[31][10] ),
    .B(_09609_),
    .Y(_09622_));
 sky130_fd_sc_hd__a211o_4 _16141_ (.A1(_09210_),
    .A2(_09617_),
    .B1(_09614_),
    .C1(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__inv_2 _16142_ (.A(_09623_),
    .Y(_00024_));
 sky130_fd_sc_hd__nor2_4 _16143_ (.A(\CPU_Xreg_value_a4[31][9] ),
    .B(_09565_),
    .Y(_09624_));
 sky130_fd_sc_hd__a211o_4 _16144_ (.A1(_09213_),
    .A2(_09617_),
    .B1(_09614_),
    .C1(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__inv_2 _16145_ (.A(_09625_),
    .Y(_00023_));
 sky130_fd_sc_hd__nor2_4 _16146_ (.A(\CPU_Xreg_value_a4[31][8] ),
    .B(_09565_),
    .Y(_09626_));
 sky130_fd_sc_hd__a211o_4 _16147_ (.A1(_09218_),
    .A2(_09617_),
    .B1(_09614_),
    .C1(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__inv_2 _16148_ (.A(_09627_),
    .Y(_00022_));
 sky130_fd_sc_hd__nor2_4 _16149_ (.A(\CPU_Xreg_value_a4[31][7] ),
    .B(_09565_),
    .Y(_09628_));
 sky130_fd_sc_hd__a211o_4 _16150_ (.A1(_09221_),
    .A2(_09617_),
    .B1(_07273_),
    .C1(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__inv_2 _16151_ (.A(_09629_),
    .Y(_00021_));
 sky130_fd_sc_hd__nor2_4 _16152_ (.A(\CPU_Xreg_value_a4[31][6] ),
    .B(_09565_),
    .Y(_09630_));
 sky130_fd_sc_hd__a211o_4 _16153_ (.A1(_09224_),
    .A2(_09569_),
    .B1(_07273_),
    .C1(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__inv_2 _16154_ (.A(_09631_),
    .Y(_00020_));
 sky130_fd_sc_hd__nor2_4 _16155_ (.A(\CPU_Xreg_value_a4[31][5] ),
    .B(_09565_),
    .Y(_09632_));
 sky130_fd_sc_hd__a211o_4 _16156_ (.A1(_09227_),
    .A2(_09569_),
    .B1(_07273_),
    .C1(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__inv_2 _16157_ (.A(_09633_),
    .Y(_00019_));
 sky130_fd_sc_hd__and2_4 _16158_ (.A(\CPU_Xreg_value_a4[31][4] ),
    .B(_09563_),
    .X(_09634_));
 sky130_fd_sc_hd__a211o_4 _16159_ (.A1(_08345_),
    .A2(_09566_),
    .B1(_09483_),
    .C1(_09634_),
    .X(_00018_));
 sky130_fd_sc_hd__and2_4 _16160_ (.A(\CPU_Xreg_value_a4[31][3] ),
    .B(_09563_),
    .X(_01550_));
 sky130_fd_sc_hd__a211o_4 _16161_ (.A1(_07641_),
    .A2(_09566_),
    .B1(_06103_),
    .C1(_01550_),
    .X(_00017_));
 sky130_fd_sc_hd__and2_4 _16162_ (.A(\CPU_Xreg_value_a4[31][2] ),
    .B(_09563_),
    .X(_01551_));
 sky130_fd_sc_hd__a211o_4 _16163_ (.A1(_07271_),
    .A2(_09566_),
    .B1(_06103_),
    .C1(_01551_),
    .X(_00016_));
 sky130_fd_sc_hd__and2_4 _16164_ (.A(\CPU_Xreg_value_a4[31][1] ),
    .B(_09563_),
    .X(_01552_));
 sky130_fd_sc_hd__a211o_4 _16165_ (.A1(_07096_),
    .A2(_09566_),
    .B1(_06103_),
    .C1(_01552_),
    .X(_00015_));
 sky130_fd_sc_hd__and2_4 _16166_ (.A(\CPU_Xreg_value_a4[31][0] ),
    .B(_09563_),
    .X(_01553_));
 sky130_fd_sc_hd__a211o_4 _16167_ (.A1(_06981_),
    .A2(_09566_),
    .B1(_06103_),
    .C1(_01553_),
    .X(_00014_));
 sky130_fd_sc_hd__inv_2 _16168_ (.A(CPU_is_blt_a3),
    .Y(_01554_));
 sky130_fd_sc_hd__inv_2 _16169_ (.A(_06934_),
    .Y(_01555_));
 sky130_fd_sc_hd__o21ai_4 _16170_ (.A1(_06493_),
    .A2(_01555_),
    .B1(_06935_),
    .Y(_01556_));
 sky130_fd_sc_hd__a32o_4 _16171_ (.A1(CPU_is_bltu_a3),
    .A2(_01554_),
    .A3(_01555_),
    .B1(CPU_is_blt_a3),
    .B2(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__buf_2 _16172_ (.A(_01557_),
    .X(_01558_));
 sky130_fd_sc_hd__inv_2 _16173_ (.A(_01557_),
    .Y(_01559_));
 sky130_fd_sc_hd__and2_4 _16174_ (.A(CPU_is_load_a3),
    .B(_06154_),
    .X(_01560_));
 sky130_fd_sc_hd__buf_2 _16175_ (.A(_01560_),
    .X(CPU_valid_load_a3));
 sky130_fd_sc_hd__inv_2 _16176_ (.A(CPU_valid_load_a3),
    .Y(_01561_));
 sky130_fd_sc_hd__buf_2 _16177_ (.A(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__o22a_4 _16178_ (.A1(\CPU_inc_pc_a1[1] ),
    .A2(CPU_valid_load_a3),
    .B1(\CPU_inc_pc_a3[1] ),
    .B2(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__a22oi_4 _16179_ (.A1(\CPU_br_tgt_pc_a3[1] ),
    .A2(_01558_),
    .B1(_01559_),
    .B2(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_4 _16180_ (.A(CPU_reset_a1),
    .B(_01564_),
    .Y(_00013_));
 sky130_fd_sc_hd__o22a_4 _16181_ (.A1(\CPU_inc_pc_a1[0] ),
    .A2(CPU_valid_load_a3),
    .B1(\CPU_inc_pc_a3[0] ),
    .B2(_01562_),
    .X(_01565_));
 sky130_fd_sc_hd__a22oi_4 _16182_ (.A1(\CPU_br_tgt_pc_a3[0] ),
    .A2(_01558_),
    .B1(_01559_),
    .B2(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_4 _16183_ (.A(CPU_reset_a1),
    .B(_01566_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _16184_ (.A(\CPU_imem_rd_addr_a1[3] ),
    .Y(_01567_));
 sky130_fd_sc_hd__buf_2 _16185_ (.A(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__buf_2 _16186_ (.A(\CPU_imem_rd_addr_a1[1] ),
    .X(_01569_));
 sky130_fd_sc_hd__and3_4 _16187_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .B(_01569_),
    .C(\CPU_imem_rd_addr_a1[2] ),
    .X(_01570_));
 sky130_fd_sc_hd__inv_2 _16188_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .Y(\CPU_inc_pc_a1[2] ));
 sky130_fd_sc_hd__inv_2 _16189_ (.A(\CPU_imem_rd_addr_a1[1] ),
    .Y(_01571_));
 sky130_fd_sc_hd__or2_4 _16190_ (.A(\CPU_inc_pc_a1[2] ),
    .B(_01571_),
    .X(_01572_));
 sky130_fd_sc_hd__inv_2 _16191_ (.A(\CPU_imem_rd_addr_a1[2] ),
    .Y(_01573_));
 sky130_fd_sc_hd__or2_4 _16192_ (.A(\CPU_imem_rd_addr_a1[3] ),
    .B(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__or2_4 _16193_ (.A(_01572_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__o21ai_4 _16194_ (.A1(_01568_),
    .A2(_01570_),
    .B1(_01575_),
    .Y(\CPU_inc_pc_a1[5] ));
 sky130_fd_sc_hd__o22a_4 _16195_ (.A1(\CPU_inc_pc_a3[5] ),
    .A2(_01562_),
    .B1(CPU_valid_load_a3),
    .B2(\CPU_inc_pc_a1[5] ),
    .X(_01576_));
 sky130_fd_sc_hd__a22oi_4 _16196_ (.A1(\CPU_br_tgt_pc_a3[5] ),
    .A2(_01558_),
    .B1(_01559_),
    .B2(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__nor2_4 _16197_ (.A(CPU_reset_a1),
    .B(_01577_),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _16198_ (.A(CPU_reset_a1),
    .Y(_01578_));
 sky130_fd_sc_hd__or2_4 _16199_ (.A(\CPU_br_tgt_pc_a3[4] ),
    .B(_01559_),
    .X(_01579_));
 sky130_fd_sc_hd__a21oi_4 _16200_ (.A1(_01573_),
    .A2(_01572_),
    .B1(_01570_),
    .Y(\CPU_inc_pc_a1[4] ));
 sky130_fd_sc_hd__and2_4 _16201_ (.A(\CPU_inc_pc_a3[4] ),
    .B(CPU_valid_load_a3),
    .X(_01580_));
 sky130_fd_sc_hd__a211o_4 _16202_ (.A1(_01562_),
    .A2(\CPU_inc_pc_a1[4] ),
    .B1(_01580_),
    .C1(_01557_),
    .X(_01581_));
 sky130_fd_sc_hd__and3_4 _16203_ (.A(_01578_),
    .B(_01579_),
    .C(_01581_),
    .X(_00010_));
 sky130_fd_sc_hd__inv_2 _16204_ (.A(\CPU_br_tgt_pc_a3[3] ),
    .Y(_01582_));
 sky130_fd_sc_hd__buf_2 _16205_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .X(_01583_));
 sky130_fd_sc_hd__o22a_4 _16206_ (.A1(\CPU_inc_pc_a1[2] ),
    .A2(_01569_),
    .B1(_01583_),
    .B2(_01571_),
    .X(_01584_));
 sky130_fd_sc_hd__a2bb2o_4 _16207_ (.A1_N(\CPU_inc_pc_a3[3] ),
    .A2_N(_01562_),
    .B1(_01562_),
    .B2(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__o22a_4 _16208_ (.A1(_01582_),
    .A2(_01559_),
    .B1(_01558_),
    .B2(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__nor2_4 _16209_ (.A(CPU_reset_a1),
    .B(_01586_),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _16210_ (.A(\CPU_br_tgt_pc_a3[2] ),
    .Y(_01587_));
 sky130_fd_sc_hd__a2bb2o_4 _16211_ (.A1_N(\CPU_inc_pc_a3[2] ),
    .A2_N(_01561_),
    .B1(_01583_),
    .B2(_01561_),
    .X(_01588_));
 sky130_fd_sc_hd__o22a_4 _16212_ (.A1(_01587_),
    .A2(_01559_),
    .B1(_01558_),
    .B2(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__nor2_4 _16213_ (.A(CPU_reset_a1),
    .B(_01589_),
    .Y(_00008_));
 sky130_fd_sc_hd__or4_4 _16214_ (.A(\CPU_Xreg_value_a5[17][21] ),
    .B(\CPU_Xreg_value_a5[17][20] ),
    .C(\CPU_Xreg_value_a5[17][23] ),
    .D(\CPU_Xreg_value_a5[17][22] ),
    .X(_01590_));
 sky130_fd_sc_hd__or4_4 _16215_ (.A(\CPU_Xreg_value_a5[17][17] ),
    .B(\CPU_Xreg_value_a5[17][16] ),
    .C(\CPU_Xreg_value_a5[17][19] ),
    .D(\CPU_Xreg_value_a5[17][18] ),
    .X(_01591_));
 sky130_fd_sc_hd__or4_4 _16216_ (.A(\CPU_Xreg_value_a5[17][29] ),
    .B(\CPU_Xreg_value_a5[17][28] ),
    .C(\CPU_Xreg_value_a5[17][31] ),
    .D(\CPU_Xreg_value_a5[17][30] ),
    .X(_01592_));
 sky130_fd_sc_hd__or4_4 _16217_ (.A(\CPU_Xreg_value_a5[17][25] ),
    .B(\CPU_Xreg_value_a5[17][24] ),
    .C(\CPU_Xreg_value_a5[17][27] ),
    .D(\CPU_Xreg_value_a5[17][26] ),
    .X(_01593_));
 sky130_fd_sc_hd__or4_4 _16218_ (.A(_01590_),
    .B(_01591_),
    .C(_01592_),
    .D(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__inv_2 _16219_ (.A(\CPU_Xreg_value_a5[17][1] ),
    .Y(_01595_));
 sky130_fd_sc_hd__and4_4 _16220_ (.A(\CPU_Xreg_value_a5[17][3] ),
    .B(\CPU_Xreg_value_a5[17][2] ),
    .C(_01595_),
    .D(\CPU_Xreg_value_a5[17][0] ),
    .X(_01596_));
 sky130_fd_sc_hd__inv_2 _16221_ (.A(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__inv_2 _16222_ (.A(\CPU_Xreg_value_a5[17][5] ),
    .Y(_01598_));
 sky130_fd_sc_hd__or4_4 _16223_ (.A(\CPU_Xreg_value_a5[17][7] ),
    .B(\CPU_Xreg_value_a5[17][6] ),
    .C(_01598_),
    .D(\CPU_Xreg_value_a5[17][4] ),
    .X(_01599_));
 sky130_fd_sc_hd__or4_4 _16224_ (.A(\CPU_Xreg_value_a5[17][13] ),
    .B(\CPU_Xreg_value_a5[17][12] ),
    .C(\CPU_Xreg_value_a5[17][15] ),
    .D(\CPU_Xreg_value_a5[17][14] ),
    .X(_01600_));
 sky130_fd_sc_hd__or4_4 _16225_ (.A(\CPU_Xreg_value_a5[17][9] ),
    .B(\CPU_Xreg_value_a5[17][8] ),
    .C(\CPU_Xreg_value_a5[17][11] ),
    .D(\CPU_Xreg_value_a5[17][10] ),
    .X(_01601_));
 sky130_fd_sc_hd__or4_4 _16226_ (.A(_01597_),
    .B(_01599_),
    .C(_01600_),
    .D(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_4 _16227_ (.A(_01594_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__and2_4 _16228_ (.A(out[7]),
    .B(_01603_),
    .X(_00007_));
 sky130_fd_sc_hd__and2_4 _16229_ (.A(out[6]),
    .B(_01603_),
    .X(_00006_));
 sky130_fd_sc_hd__inv_2 _16230_ (.A(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__or2_4 _16231_ (.A(out[5]),
    .B(_01604_),
    .X(_00005_));
 sky130_fd_sc_hd__and2_4 _16232_ (.A(out[4]),
    .B(_01603_),
    .X(_00004_));
 sky130_fd_sc_hd__or2_4 _16233_ (.A(out[3]),
    .B(_01604_),
    .X(_00003_));
 sky130_fd_sc_hd__or2_4 _16234_ (.A(out[2]),
    .B(_01604_),
    .X(_00002_));
 sky130_fd_sc_hd__and2_4 _16235_ (.A(out[1]),
    .B(_01603_),
    .X(_00001_));
 sky130_fd_sc_hd__or2_4 _16236_ (.A(out[0]),
    .B(_01604_),
    .X(_00000_));
 sky130_fd_sc_hd__or3_4 _16237_ (.A(\CPU_imem_rd_addr_a1[1] ),
    .B(_01567_),
    .C(\CPU_imem_rd_addr_a1[2] ),
    .X(_01605_));
 sky130_fd_sc_hd__buf_2 _16238_ (.A(_01605_),
    .X(\CPU_imem_rd_data_a1[10] ));
 sky130_fd_sc_hd__inv_2 _16239_ (.A(\CPU_imem_rd_data_a1[10] ),
    .Y(_01606_));
 sky130_fd_sc_hd__and2_4 _16240_ (.A(\CPU_inc_pc_a1[2] ),
    .B(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_2 _16241_ (.A(_01607_),
    .X(CPU_is_s_instr_a1));
 sky130_fd_sc_hd__inv_2 _16242_ (.A(_01574_),
    .Y(\CPU_imem_rd_data_a1[17] ));
 sky130_fd_sc_hd__and2_4 _16243_ (.A(\CPU_inc_pc_a1[2] ),
    .B(\CPU_imem_rd_data_a1[17] ),
    .X(_01608_));
 sky130_fd_sc_hd__buf_2 _16244_ (.A(_01608_),
    .X(\CPU_imem_rd_data_a1[22] ));
 sky130_fd_sc_hd__and2_4 _16245_ (.A(_01569_),
    .B(\CPU_imem_rd_data_a1[22] ),
    .X(_01609_));
 sky130_fd_sc_hd__buf_2 _16246_ (.A(_01609_),
    .X(CPU_is_blt_a1));
 sky130_fd_sc_hd__and2_4 _16247_ (.A(_01606_),
    .B(CPU_is_blt_a1),
    .X(CPU_is_bltu_a1));
 sky130_fd_sc_hd__and4_4 _16248_ (.A(_01583_),
    .B(_01571_),
    .C(_01568_),
    .D(_01573_),
    .X(_01610_));
 sky130_fd_sc_hd__or2_4 _16249_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .B(\CPU_imem_rd_addr_a1[1] ),
    .X(_01611_));
 sky130_fd_sc_hd__and3_4 _16250_ (.A(_01567_),
    .B(_01573_),
    .C(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__or2_4 _16251_ (.A(\CPU_imem_rd_data_a1[17] ),
    .B(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__nor2_4 _16252_ (.A(_01606_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__or4_4 _16253_ (.A(_01584_),
    .B(_01610_),
    .C(CPU_is_blt_a1),
    .D(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__inv_2 _16254_ (.A(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__or2_4 _16255_ (.A(CPU_is_s_instr_a1),
    .B(_01609_),
    .X(_01617_));
 sky130_fd_sc_hd__and2_4 _16256_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .B(_01606_),
    .X(_01618_));
 sky130_fd_sc_hd__buf_2 _16257_ (.A(_01618_),
    .X(CPU_is_load_a1));
 sky130_fd_sc_hd__or2_4 _16258_ (.A(_01617_),
    .B(CPU_is_load_a1),
    .X(_01619_));
 sky130_fd_sc_hd__buf_2 _16259_ (.A(_01619_),
    .X(\CPU_imem_rd_data_a1[11] ));
 sky130_fd_sc_hd__nor2_4 _16260_ (.A(_01616_),
    .B(\CPU_imem_rd_data_a1[11] ),
    .Y(CPU_is_add_a1));
 sky130_fd_sc_hd__nor2_4 _16261_ (.A(_01615_),
    .B(\CPU_imem_rd_data_a1[11] ),
    .Y(CPU_is_addi_a1));
 sky130_fd_sc_hd__inv_2 _16262_ (.A(_01617_),
    .Y(\gen_clkP_CPU_rd_valid_a2.pwr_en ));
 sky130_fd_sc_hd__and2_4 _16263_ (.A(CPU_valid_a3),
    .B(_01558_),
    .X(CPU_valid_taken_br_a3));
 sky130_fd_sc_hd__and4_4 _16264_ (.A(_01583_),
    .B(_01569_),
    .C(_01568_),
    .D(_01573_),
    .X(_01620_));
 sky130_fd_sc_hd__and4_4 _16265_ (.A(_01568_),
    .B(\CPU_imem_rd_addr_a1[2] ),
    .C(_01571_),
    .D(_01583_),
    .X(_01621_));
 sky130_fd_sc_hd__buf_2 _16266_ (.A(_01621_),
    .X(\CPU_imem_rd_data_a1[20] ));
 sky130_fd_sc_hd__or4_4 _16267_ (.A(CPU_is_blt_a1),
    .B(_01620_),
    .C(CPU_is_load_a1),
    .D(\CPU_imem_rd_data_a1[20] ),
    .X(\CPU_imem_rd_data_a1[7] ));
 sky130_fd_sc_hd__inv_2 _16268_ (.A(_01575_),
    .Y(_01622_));
 sky130_fd_sc_hd__and2_4 _16269_ (.A(_01571_),
    .B(\CPU_imem_rd_data_a1[22] ),
    .X(_01623_));
 sky130_fd_sc_hd__or4_4 _16270_ (.A(_01622_),
    .B(_01610_),
    .C(_01623_),
    .D(_01614_),
    .X(\CPU_imem_rd_data_a1[8] ));
 sky130_fd_sc_hd__a21o_4 _16271_ (.A1(_01571_),
    .A2(\CPU_imem_rd_data_a1[17] ),
    .B1(_01612_),
    .X(\CPU_imem_rd_data_a1[9] ));
 sky130_fd_sc_hd__and2_4 _16272_ (.A(_01572_),
    .B(\CPU_imem_rd_data_a1[17] ),
    .X(\CPU_imem_rd_data_a1[15] ));
 sky130_fd_sc_hd__or2_4 _16273_ (.A(_01622_),
    .B(_01612_),
    .X(\CPU_imem_rd_data_a1[16] ));
 sky130_fd_sc_hd__and2_4 _16274_ (.A(_01568_),
    .B(_01613_),
    .X(\CPU_imem_rd_data_a1[18] ));
 sky130_fd_sc_hd__and4_4 _16275_ (.A(\CPU_inc_pc_a1[2] ),
    .B(_01569_),
    .C(_01568_),
    .D(_01573_),
    .X(\CPU_imm_a1[1] ));
 sky130_fd_sc_hd__or3_4 _16276_ (.A(CPU_is_s_instr_a1),
    .B(\CPU_imm_a1[1] ),
    .C(_01623_),
    .X(\CPU_imem_rd_data_a1[21] ));
 sky130_fd_sc_hd__nor2_4 _16277_ (.A(_01583_),
    .B(_01614_),
    .Y(\CPU_imem_rd_data_a1[23] ));
 sky130_fd_sc_hd__buf_2 _16278_ (.A(CPU_is_load_a1),
    .X(\CPU_imem_rd_data_a1[24] ));
 sky130_fd_sc_hd__inv_2 _16279_ (.A(_01584_),
    .Y(\CPU_inc_pc_a1[3] ));
 sky130_fd_sc_hd__buf_2 _16280_ (.A(\CPU_imem_rd_data_a1[20] ),
    .X(\CPU_imm_a1[0] ));
 sky130_fd_sc_hd__and2_4 _16281_ (.A(\CPU_imem_rd_data_a1[22] ),
    .B(_01616_),
    .X(\CPU_imm_a1[2] ));
 sky130_fd_sc_hd__and2_4 _16282_ (.A(_01569_),
    .B(\CPU_imem_rd_data_a1[23] ),
    .X(\CPU_imm_a1[3] ));
 sky130_fd_sc_hd__buf_2 _16283_ (.A(\CPU_imem_rd_data_a1[11] ),
    .X(\CPU_imm_a1[4] ));
 sky130_fd_sc_hd__buf_2 _16284_ (.A(CPU_is_blt_a1),
    .X(\CPU_imm_a1[10] ));
 sky130_fd_sc_hd__buf_2 _16285_ (.A(CPU_is_blt_a1),
    .X(\CPU_imm_a1[11] ));
 sky130_fd_sc_hd__inv_2 _16286_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .Y(_01624_));
 sky130_fd_sc_hd__buf_2 _16287_ (.A(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_4 _16288_ (.A(\CPU_rd_a3[1] ),
    .B(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__inv_2 _16289_ (.A(\CPU_rf_rd_index1_a2[3] ),
    .Y(_01627_));
 sky130_fd_sc_hd__buf_2 _16290_ (.A(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__a2bb2o_4 _16291_ (.A1_N(\CPU_rd_a3[1] ),
    .A2_N(_01625_),
    .B1(\CPU_rd_a3[3] ),
    .B2(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__inv_2 _16292_ (.A(\CPU_rd_a3[2] ),
    .Y(_01630_));
 sky130_fd_sc_hd__buf_2 _16293_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .X(_01631_));
 sky130_fd_sc_hd__and2_4 _16294_ (.A(_01630_),
    .B(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__inv_2 _16295_ (.A(\CPU_rd_a3[3] ),
    .Y(_01633_));
 sky130_fd_sc_hd__buf_2 _16296_ (.A(\CPU_rf_rd_index1_a2[3] ),
    .X(_01634_));
 sky130_fd_sc_hd__a2bb2o_4 _16297_ (.A1_N(_01630_),
    .A2_N(_01631_),
    .B1(_01633_),
    .B2(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__buf_2 _16298_ (.A(\CPU_rf_rd_index1_a2[0] ),
    .X(_01636_));
 sky130_fd_sc_hd__inv_2 _16299_ (.A(\CPU_rd_a3[0] ),
    .Y(_01637_));
 sky130_fd_sc_hd__inv_2 _16300_ (.A(\CPU_rf_rd_index1_a2[0] ),
    .Y(_01638_));
 sky130_fd_sc_hd__buf_2 _16301_ (.A(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__o22a_4 _16302_ (.A1(\CPU_rd_a3[0] ),
    .A2(_01636_),
    .B1(_01637_),
    .B2(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__or4_4 _16303_ (.A(\CPU_rd_a3[4] ),
    .B(_01632_),
    .C(_01635_),
    .D(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__inv_2 _16304_ (.A(_06162_),
    .Y(_01642_));
 sky130_fd_sc_hd__or4_4 _16305_ (.A(_01626_),
    .B(_01629_),
    .C(_01641_),
    .D(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__buf_2 _16306_ (.A(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__buf_2 _16307_ (.A(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__inv_2 _16308_ (.A(_01643_),
    .Y(_01646_));
 sky130_fd_sc_hd__buf_2 _16309_ (.A(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__buf_2 _16310_ (.A(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__or4_4 _16311_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .C(\CPU_rf_rd_index1_a2[2] ),
    .D(\CPU_rf_rd_index1_a2[3] ),
    .X(_01649_));
 sky130_fd_sc_hd__buf_2 _16312_ (.A(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__buf_2 _16313_ (.A(_01650_),
    .X(_01651_));
 sky130_fd_sc_hd__buf_2 _16314_ (.A(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__buf_2 _16315_ (.A(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__inv_2 _16316_ (.A(\CPU_Xreg_value_a4[8][0] ),
    .Y(_01654_));
 sky130_fd_sc_hd__buf_2 _16317_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .X(_01655_));
 sky130_fd_sc_hd__or4_4 _16318_ (.A(_01655_),
    .B(_01636_),
    .C(_01631_),
    .D(_01628_),
    .X(_01656_));
 sky130_fd_sc_hd__buf_2 _16319_ (.A(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__inv_2 _16320_ (.A(\CPU_Xreg_value_a4[13][0] ),
    .Y(_01658_));
 sky130_fd_sc_hd__inv_2 _16321_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .Y(_01659_));
 sky130_fd_sc_hd__buf_2 _16322_ (.A(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__or4_4 _16323_ (.A(_01660_),
    .B(_01628_),
    .C(_01655_),
    .D(_01639_),
    .X(_01661_));
 sky130_fd_sc_hd__o22a_4 _16324_ (.A1(_01654_),
    .A2(_01657_),
    .B1(_01658_),
    .B2(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__or4_4 _16325_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(_01638_),
    .C(_01659_),
    .D(\CPU_rf_rd_index1_a2[3] ),
    .X(_01663_));
 sky130_fd_sc_hd__buf_2 _16326_ (.A(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__buf_2 _16327_ (.A(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__inv_2 _16328_ (.A(\CPU_Xreg_value_a4[12][0] ),
    .Y(_01666_));
 sky130_fd_sc_hd__or4_4 _16329_ (.A(_01655_),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .C(_01659_),
    .D(_01627_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_2 _16330_ (.A(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__buf_2 _16331_ (.A(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__o22a_4 _16332_ (.A1(_07363_),
    .A2(_01665_),
    .B1(_01666_),
    .B2(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__inv_2 _16333_ (.A(\CPU_Xreg_value_a4[2][0] ),
    .Y(_01671_));
 sky130_fd_sc_hd__or4_4 _16334_ (.A(_01631_),
    .B(_01634_),
    .C(_01625_),
    .D(_01636_),
    .X(_01672_));
 sky130_fd_sc_hd__buf_2 _16335_ (.A(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__o21a_4 _16336_ (.A1(_01671_),
    .A2(_01673_),
    .B1(_01651_),
    .X(_01674_));
 sky130_fd_sc_hd__inv_2 _16337_ (.A(\CPU_Xreg_value_a4[14][0] ),
    .Y(_01675_));
 sky130_fd_sc_hd__or4_4 _16338_ (.A(_01660_),
    .B(_01627_),
    .C(_01624_),
    .D(\CPU_rf_rd_index1_a2[0] ),
    .X(_01676_));
 sky130_fd_sc_hd__buf_2 _16339_ (.A(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__buf_2 _16340_ (.A(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__or4_4 _16341_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .C(_01624_),
    .D(_01638_),
    .X(_01679_));
 sky130_fd_sc_hd__buf_2 _16342_ (.A(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__buf_2 _16343_ (.A(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__o22a_4 _16344_ (.A1(_01675_),
    .A2(_01678_),
    .B1(_07189_),
    .B2(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__and4_4 _16345_ (.A(_01662_),
    .B(_01670_),
    .C(_01674_),
    .D(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__or4_4 _16346_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(_01634_),
    .C(_01655_),
    .D(_01639_),
    .X(_01684_));
 sky130_fd_sc_hd__buf_2 _16347_ (.A(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__buf_2 _16348_ (.A(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__inv_2 _16349_ (.A(\CPU_Xreg_value_a4[4][0] ),
    .Y(_01687_));
 sky130_fd_sc_hd__or4_4 _16350_ (.A(_01655_),
    .B(_01636_),
    .C(_01660_),
    .D(_01634_),
    .X(_01688_));
 sky130_fd_sc_hd__buf_2 _16351_ (.A(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__buf_2 _16352_ (.A(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__o22a_4 _16353_ (.A1(_06982_),
    .A2(_01686_),
    .B1(_01687_),
    .B2(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__inv_2 _16354_ (.A(\CPU_Xreg_value_a4[6][0] ),
    .Y(_01692_));
 sky130_fd_sc_hd__or4_4 _16355_ (.A(_01660_),
    .B(_01634_),
    .C(_01624_),
    .D(_01636_),
    .X(_01693_));
 sky130_fd_sc_hd__buf_2 _16356_ (.A(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__buf_2 _16357_ (.A(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__or4_4 _16358_ (.A(_01631_),
    .B(_01628_),
    .C(_01625_),
    .D(_01639_),
    .X(_01696_));
 sky130_fd_sc_hd__buf_2 _16359_ (.A(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__buf_2 _16360_ (.A(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__o22a_4 _16361_ (.A1(_01692_),
    .A2(_01695_),
    .B1(_07902_),
    .B2(_01698_),
    .X(_01699_));
 sky130_fd_sc_hd__or4_4 _16362_ (.A(_01660_),
    .B(_01628_),
    .C(_01624_),
    .D(_01639_),
    .X(_01700_));
 sky130_fd_sc_hd__buf_2 _16363_ (.A(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__buf_2 _16364_ (.A(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__inv_2 _16365_ (.A(\CPU_Xreg_value_a4[10][0] ),
    .Y(_01703_));
 sky130_fd_sc_hd__or4_4 _16366_ (.A(_01631_),
    .B(_01628_),
    .C(_01625_),
    .D(_01636_),
    .X(_01704_));
 sky130_fd_sc_hd__buf_2 _16367_ (.A(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__buf_2 _16368_ (.A(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__o22a_4 _16369_ (.A1(_08271_),
    .A2(_01702_),
    .B1(_01703_),
    .B2(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__or4_4 _16370_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(_01627_),
    .C(_01655_),
    .D(_01638_),
    .X(_01708_));
 sky130_fd_sc_hd__buf_2 _16371_ (.A(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__buf_2 _16372_ (.A(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__or4_4 _16373_ (.A(_01660_),
    .B(_01634_),
    .C(_01625_),
    .D(_01639_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_2 _16374_ (.A(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__buf_2 _16375_ (.A(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__o22a_4 _16376_ (.A1(_07733_),
    .A2(_01710_),
    .B1(_07533_),
    .B2(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__and4_4 _16377_ (.A(_01691_),
    .B(_01699_),
    .C(_01707_),
    .D(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__a2bb2o_4 _16378_ (.A1_N(\CPU_Xreg_value_a4[0][0] ),
    .A2_N(_01653_),
    .B1(_01683_),
    .B2(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__inv_2 _16379_ (.A(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__o22a_4 _16380_ (.A1(_06979_),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01717_),
    .X(\CPU_src1_value_a2[0] ));
 sky130_fd_sc_hd__buf_2 _16381_ (.A(_01653_),
    .X(_01718_));
 sky130_fd_sc_hd__inv_2 _16382_ (.A(\CPU_Xreg_value_a4[8][1] ),
    .Y(_01719_));
 sky130_fd_sc_hd__buf_2 _16383_ (.A(_01657_),
    .X(_01720_));
 sky130_fd_sc_hd__inv_2 _16384_ (.A(_01661_),
    .Y(_01721_));
 sky130_fd_sc_hd__buf_2 _16385_ (.A(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__a2bb2o_4 _16386_ (.A1_N(_01719_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][1] ),
    .B2(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__inv_2 _16387_ (.A(\CPU_Xreg_value_a4[5][1] ),
    .Y(_01724_));
 sky130_fd_sc_hd__inv_2 _16388_ (.A(\CPU_Xreg_value_a4[12][1] ),
    .Y(_01725_));
 sky130_fd_sc_hd__o22a_4 _16389_ (.A1(_01724_),
    .A2(_01665_),
    .B1(_01725_),
    .B2(_01669_),
    .X(_01726_));
 sky130_fd_sc_hd__inv_2 _16390_ (.A(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__buf_2 _16391_ (.A(_01673_),
    .X(_01728_));
 sky130_fd_sc_hd__o21ai_4 _16392_ (.A1(_07098_),
    .A2(_01728_),
    .B1(_01652_),
    .Y(_01729_));
 sky130_fd_sc_hd__o22a_4 _16393_ (.A1(_08182_),
    .A2(_01678_),
    .B1(_07186_),
    .B2(_01681_),
    .X(_01730_));
 sky130_fd_sc_hd__inv_2 _16394_ (.A(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__or4_4 _16395_ (.A(_01723_),
    .B(_01727_),
    .C(_01729_),
    .D(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__inv_2 _16396_ (.A(\CPU_Xreg_value_a4[1][1] ),
    .Y(_01733_));
 sky130_fd_sc_hd__inv_2 _16397_ (.A(\CPU_Xreg_value_a4[4][1] ),
    .Y(_01734_));
 sky130_fd_sc_hd__o22a_4 _16398_ (.A1(_01733_),
    .A2(_01686_),
    .B1(_01734_),
    .B2(_01690_),
    .X(_01735_));
 sky130_fd_sc_hd__o22a_4 _16399_ (.A1(_07445_),
    .A2(_01695_),
    .B1(_07900_),
    .B2(_01698_),
    .X(_01736_));
 sky130_fd_sc_hd__o22a_4 _16400_ (.A1(_08268_),
    .A2(_01702_),
    .B1(_07817_),
    .B2(_01706_),
    .X(_01737_));
 sky130_fd_sc_hd__inv_2 _16401_ (.A(\CPU_Xreg_value_a4[9][1] ),
    .Y(_01738_));
 sky130_fd_sc_hd__o22a_4 _16402_ (.A1(_01738_),
    .A2(_01710_),
    .B1(_07531_),
    .B2(_01713_),
    .X(_01739_));
 sky130_fd_sc_hd__and4_4 _16403_ (.A(_01735_),
    .B(_01736_),
    .C(_01737_),
    .D(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__inv_2 _16404_ (.A(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__o22a_4 _16405_ (.A1(\CPU_Xreg_value_a4[0][1] ),
    .A2(_01718_),
    .B1(_01732_),
    .B2(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__o22a_4 _16406_ (.A1(_06866_),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01742_),
    .X(\CPU_src1_value_a2[1] ));
 sky130_fd_sc_hd__inv_2 _16407_ (.A(\CPU_Xreg_value_a4[8][2] ),
    .Y(_01743_));
 sky130_fd_sc_hd__a2bb2o_4 _16408_ (.A1_N(_01743_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][2] ),
    .B2(_01722_),
    .X(_01744_));
 sky130_fd_sc_hd__o22a_4 _16409_ (.A1(_07359_),
    .A2(_01665_),
    .B1(_07983_),
    .B2(_01669_),
    .X(_01745_));
 sky130_fd_sc_hd__inv_2 _16410_ (.A(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__inv_2 _16411_ (.A(\CPU_Xreg_value_a4[2][2] ),
    .Y(_01747_));
 sky130_fd_sc_hd__o21ai_4 _16412_ (.A1(_01747_),
    .A2(_01728_),
    .B1(_01652_),
    .Y(_01748_));
 sky130_fd_sc_hd__inv_2 _16413_ (.A(\CPU_Xreg_value_a4[3][2] ),
    .Y(_01749_));
 sky130_fd_sc_hd__o22a_4 _16414_ (.A1(_08179_),
    .A2(_01678_),
    .B1(_01749_),
    .B2(_01681_),
    .X(_01750_));
 sky130_fd_sc_hd__inv_2 _16415_ (.A(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__or4_4 _16416_ (.A(_01744_),
    .B(_01746_),
    .C(_01748_),
    .D(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__inv_2 _16417_ (.A(\CPU_Xreg_value_a4[1][2] ),
    .Y(_01753_));
 sky130_fd_sc_hd__o22a_4 _16418_ (.A1(_01753_),
    .A2(_01686_),
    .B1(_07275_),
    .B2(_01690_),
    .X(_01754_));
 sky130_fd_sc_hd__inv_2 _16419_ (.A(\CPU_Xreg_value_a4[11][2] ),
    .Y(_01755_));
 sky130_fd_sc_hd__o22a_4 _16420_ (.A1(_07443_),
    .A2(_01695_),
    .B1(_01755_),
    .B2(_01698_),
    .X(_01756_));
 sky130_fd_sc_hd__inv_2 _16421_ (.A(\CPU_Xreg_value_a4[10][2] ),
    .Y(_01757_));
 sky130_fd_sc_hd__o22a_4 _16422_ (.A1(_08266_),
    .A2(_01702_),
    .B1(_01757_),
    .B2(_01706_),
    .X(_01758_));
 sky130_fd_sc_hd__inv_2 _16423_ (.A(\CPU_Xreg_value_a4[9][2] ),
    .Y(_01759_));
 sky130_fd_sc_hd__o22a_4 _16424_ (.A1(_01759_),
    .A2(_01710_),
    .B1(_07528_),
    .B2(_01713_),
    .X(_01760_));
 sky130_fd_sc_hd__and4_4 _16425_ (.A(_01754_),
    .B(_01756_),
    .C(_01758_),
    .D(_01760_),
    .X(_01761_));
 sky130_fd_sc_hd__inv_2 _16426_ (.A(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__o22a_4 _16427_ (.A1(\CPU_Xreg_value_a4[0][2] ),
    .A2(_01718_),
    .B1(_01752_),
    .B2(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__o22a_4 _16428_ (.A1(\CPU_result_a3[2] ),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01763_),
    .X(\CPU_src1_value_a2[2] ));
 sky130_fd_sc_hd__a2bb2o_4 _16429_ (.A1_N(_07643_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][3] ),
    .B2(_01722_),
    .X(_01764_));
 sky130_fd_sc_hd__inv_2 _16430_ (.A(\CPU_Xreg_value_a4[5][3] ),
    .Y(_01765_));
 sky130_fd_sc_hd__o22a_4 _16431_ (.A1(_01765_),
    .A2(_01665_),
    .B1(_07981_),
    .B2(_01669_),
    .X(_01766_));
 sky130_fd_sc_hd__inv_2 _16432_ (.A(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _16433_ (.A(\CPU_Xreg_value_a4[2][3] ),
    .Y(_01768_));
 sky130_fd_sc_hd__o21ai_4 _16434_ (.A1(_01768_),
    .A2(_01728_),
    .B1(_01652_),
    .Y(_01769_));
 sky130_fd_sc_hd__inv_2 _16435_ (.A(\CPU_Xreg_value_a4[3][3] ),
    .Y(_01770_));
 sky130_fd_sc_hd__o22a_4 _16436_ (.A1(_08176_),
    .A2(_01678_),
    .B1(_01770_),
    .B2(_01681_),
    .X(_01771_));
 sky130_fd_sc_hd__inv_2 _16437_ (.A(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__or4_4 _16438_ (.A(_01764_),
    .B(_01767_),
    .C(_01769_),
    .D(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__inv_2 _16439_ (.A(\CPU_Xreg_value_a4[1][3] ),
    .Y(_01774_));
 sky130_fd_sc_hd__inv_2 _16440_ (.A(\CPU_Xreg_value_a4[4][3] ),
    .Y(_01775_));
 sky130_fd_sc_hd__o22a_4 _16441_ (.A1(_01774_),
    .A2(_01686_),
    .B1(_01775_),
    .B2(_01690_),
    .X(_01776_));
 sky130_fd_sc_hd__inv_2 _16442_ (.A(\CPU_Xreg_value_a4[6][3] ),
    .Y(_01777_));
 sky130_fd_sc_hd__o22a_4 _16443_ (.A1(_01777_),
    .A2(_01695_),
    .B1(_07896_),
    .B2(_01698_),
    .X(_01778_));
 sky130_fd_sc_hd__o22a_4 _16444_ (.A1(_08264_),
    .A2(_01702_),
    .B1(_07812_),
    .B2(_01706_),
    .X(_01779_));
 sky130_fd_sc_hd__inv_2 _16445_ (.A(\CPU_Xreg_value_a4[7][3] ),
    .Y(_01780_));
 sky130_fd_sc_hd__o22a_4 _16446_ (.A1(_07727_),
    .A2(_01710_),
    .B1(_01780_),
    .B2(_01713_),
    .X(_01781_));
 sky130_fd_sc_hd__and4_4 _16447_ (.A(_01776_),
    .B(_01778_),
    .C(_01779_),
    .D(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__inv_2 _16448_ (.A(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__o22a_4 _16449_ (.A1(\CPU_Xreg_value_a4[0][3] ),
    .A2(_01718_),
    .B1(_01773_),
    .B2(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__o22a_4 _16450_ (.A1(\CPU_result_a3[3] ),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01784_),
    .X(\CPU_src1_value_a2[3] ));
 sky130_fd_sc_hd__inv_2 _16451_ (.A(\CPU_Xreg_value_a4[8][4] ),
    .Y(_01785_));
 sky130_fd_sc_hd__a2bb2o_4 _16452_ (.A1_N(_01785_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][4] ),
    .B2(_01722_),
    .X(_01786_));
 sky130_fd_sc_hd__inv_2 _16453_ (.A(\CPU_Xreg_value_a4[5][4] ),
    .Y(_01787_));
 sky130_fd_sc_hd__inv_2 _16454_ (.A(\CPU_Xreg_value_a4[12][4] ),
    .Y(_01788_));
 sky130_fd_sc_hd__o22a_4 _16455_ (.A1(_01787_),
    .A2(_01665_),
    .B1(_01788_),
    .B2(_01669_),
    .X(_01789_));
 sky130_fd_sc_hd__inv_2 _16456_ (.A(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__inv_2 _16457_ (.A(\CPU_Xreg_value_a4[2][4] ),
    .Y(_01791_));
 sky130_fd_sc_hd__o21ai_4 _16458_ (.A1(_01791_),
    .A2(_01728_),
    .B1(_01652_),
    .Y(_01792_));
 sky130_fd_sc_hd__inv_2 _16459_ (.A(\CPU_Xreg_value_a4[14][4] ),
    .Y(_01793_));
 sky130_fd_sc_hd__inv_2 _16460_ (.A(\CPU_Xreg_value_a4[3][4] ),
    .Y(_01794_));
 sky130_fd_sc_hd__o22a_4 _16461_ (.A1(_01793_),
    .A2(_01678_),
    .B1(_01794_),
    .B2(_01681_),
    .X(_01795_));
 sky130_fd_sc_hd__inv_2 _16462_ (.A(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__or4_4 _16463_ (.A(_01786_),
    .B(_01790_),
    .C(_01792_),
    .D(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__inv_2 _16464_ (.A(\CPU_Xreg_value_a4[1][4] ),
    .Y(_01798_));
 sky130_fd_sc_hd__inv_2 _16465_ (.A(\CPU_Xreg_value_a4[4][4] ),
    .Y(_01799_));
 sky130_fd_sc_hd__o22a_4 _16466_ (.A1(_01798_),
    .A2(_01686_),
    .B1(_01799_),
    .B2(_01690_),
    .X(_01800_));
 sky130_fd_sc_hd__inv_2 _16467_ (.A(\CPU_Xreg_value_a4[6][4] ),
    .Y(_01801_));
 sky130_fd_sc_hd__inv_2 _16468_ (.A(\CPU_Xreg_value_a4[11][4] ),
    .Y(_01802_));
 sky130_fd_sc_hd__o22a_4 _16469_ (.A1(_01801_),
    .A2(_01695_),
    .B1(_01802_),
    .B2(_01698_),
    .X(_01803_));
 sky130_fd_sc_hd__inv_2 _16470_ (.A(\CPU_Xreg_value_a4[15][4] ),
    .Y(_01804_));
 sky130_fd_sc_hd__inv_2 _16471_ (.A(\CPU_Xreg_value_a4[10][4] ),
    .Y(_01805_));
 sky130_fd_sc_hd__o22a_4 _16472_ (.A1(_01804_),
    .A2(_01702_),
    .B1(_01805_),
    .B2(_01706_),
    .X(_01806_));
 sky130_fd_sc_hd__inv_2 _16473_ (.A(\CPU_Xreg_value_a4[9][4] ),
    .Y(_01807_));
 sky130_fd_sc_hd__inv_2 _16474_ (.A(\CPU_Xreg_value_a4[7][4] ),
    .Y(_01808_));
 sky130_fd_sc_hd__o22a_4 _16475_ (.A1(_01807_),
    .A2(_01710_),
    .B1(_01808_),
    .B2(_01713_),
    .X(_01809_));
 sky130_fd_sc_hd__and4_4 _16476_ (.A(_01800_),
    .B(_01803_),
    .C(_01806_),
    .D(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__inv_2 _16477_ (.A(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__o22a_4 _16478_ (.A1(\CPU_Xreg_value_a4[0][4] ),
    .A2(_01718_),
    .B1(_01797_),
    .B2(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__o22a_4 _16479_ (.A1(\CPU_result_a3[4] ),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01812_),
    .X(\CPU_src1_value_a2[4] ));
 sky130_fd_sc_hd__inv_2 _16480_ (.A(\CPU_Xreg_value_a4[8][5] ),
    .Y(_01813_));
 sky130_fd_sc_hd__a2bb2o_4 _16481_ (.A1_N(_01813_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][5] ),
    .B2(_01722_),
    .X(_01814_));
 sky130_fd_sc_hd__inv_2 _16482_ (.A(\CPU_Xreg_value_a4[5][5] ),
    .Y(_01815_));
 sky130_fd_sc_hd__inv_2 _16483_ (.A(\CPU_Xreg_value_a4[12][5] ),
    .Y(_01816_));
 sky130_fd_sc_hd__o22a_4 _16484_ (.A1(_01815_),
    .A2(_01665_),
    .B1(_01816_),
    .B2(_01669_),
    .X(_01817_));
 sky130_fd_sc_hd__inv_2 _16485_ (.A(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _16486_ (.A(\CPU_Xreg_value_a4[2][5] ),
    .Y(_01819_));
 sky130_fd_sc_hd__buf_2 _16487_ (.A(_01651_),
    .X(_01820_));
 sky130_fd_sc_hd__o21ai_4 _16488_ (.A1(_01819_),
    .A2(_01728_),
    .B1(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__inv_2 _16489_ (.A(\CPU_Xreg_value_a4[14][5] ),
    .Y(_01822_));
 sky130_fd_sc_hd__inv_2 _16490_ (.A(\CPU_Xreg_value_a4[3][5] ),
    .Y(_01823_));
 sky130_fd_sc_hd__o22a_4 _16491_ (.A1(_01822_),
    .A2(_01678_),
    .B1(_01823_),
    .B2(_01681_),
    .X(_01824_));
 sky130_fd_sc_hd__inv_2 _16492_ (.A(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__or4_4 _16493_ (.A(_01814_),
    .B(_01818_),
    .C(_01821_),
    .D(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__inv_2 _16494_ (.A(\CPU_Xreg_value_a4[1][5] ),
    .Y(_01827_));
 sky130_fd_sc_hd__inv_2 _16495_ (.A(\CPU_Xreg_value_a4[4][5] ),
    .Y(_01828_));
 sky130_fd_sc_hd__o22a_4 _16496_ (.A1(_01827_),
    .A2(_01686_),
    .B1(_01828_),
    .B2(_01690_),
    .X(_01829_));
 sky130_fd_sc_hd__inv_2 _16497_ (.A(\CPU_Xreg_value_a4[6][5] ),
    .Y(_01830_));
 sky130_fd_sc_hd__inv_2 _16498_ (.A(\CPU_Xreg_value_a4[11][5] ),
    .Y(_01831_));
 sky130_fd_sc_hd__o22a_4 _16499_ (.A1(_01830_),
    .A2(_01695_),
    .B1(_01831_),
    .B2(_01698_),
    .X(_01832_));
 sky130_fd_sc_hd__inv_2 _16500_ (.A(\CPU_Xreg_value_a4[15][5] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _16501_ (.A(\CPU_Xreg_value_a4[10][5] ),
    .Y(_01834_));
 sky130_fd_sc_hd__o22a_4 _16502_ (.A1(_01833_),
    .A2(_01702_),
    .B1(_01834_),
    .B2(_01706_),
    .X(_01835_));
 sky130_fd_sc_hd__inv_2 _16503_ (.A(\CPU_Xreg_value_a4[9][5] ),
    .Y(_01836_));
 sky130_fd_sc_hd__inv_2 _16504_ (.A(\CPU_Xreg_value_a4[7][5] ),
    .Y(_01837_));
 sky130_fd_sc_hd__o22a_4 _16505_ (.A1(_01836_),
    .A2(_01710_),
    .B1(_01837_),
    .B2(_01713_),
    .X(_01838_));
 sky130_fd_sc_hd__and4_4 _16506_ (.A(_01829_),
    .B(_01832_),
    .C(_01835_),
    .D(_01838_),
    .X(_01839_));
 sky130_fd_sc_hd__inv_2 _16507_ (.A(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__o22a_4 _16508_ (.A1(\CPU_Xreg_value_a4[0][5] ),
    .A2(_01718_),
    .B1(_01826_),
    .B2(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__o22a_4 _16509_ (.A1(\CPU_result_a3[5] ),
    .A2(_01645_),
    .B1(_01648_),
    .B2(_01841_),
    .X(\CPU_src1_value_a2[5] ));
 sky130_fd_sc_hd__buf_2 _16510_ (.A(_01644_),
    .X(_01842_));
 sky130_fd_sc_hd__buf_2 _16511_ (.A(_01647_),
    .X(_01843_));
 sky130_fd_sc_hd__inv_2 _16512_ (.A(\CPU_Xreg_value_a4[8][6] ),
    .Y(_01844_));
 sky130_fd_sc_hd__a2bb2o_4 _16513_ (.A1_N(_01844_),
    .A2_N(_01720_),
    .B1(\CPU_Xreg_value_a4[13][6] ),
    .B2(_01722_),
    .X(_01845_));
 sky130_fd_sc_hd__inv_2 _16514_ (.A(\CPU_Xreg_value_a4[5][6] ),
    .Y(_01846_));
 sky130_fd_sc_hd__buf_2 _16515_ (.A(_01664_),
    .X(_01847_));
 sky130_fd_sc_hd__inv_2 _16516_ (.A(\CPU_Xreg_value_a4[12][6] ),
    .Y(_01848_));
 sky130_fd_sc_hd__buf_2 _16517_ (.A(_01668_),
    .X(_01849_));
 sky130_fd_sc_hd__o22a_4 _16518_ (.A1(_01846_),
    .A2(_01847_),
    .B1(_01848_),
    .B2(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__inv_2 _16519_ (.A(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__inv_2 _16520_ (.A(\CPU_Xreg_value_a4[2][6] ),
    .Y(_01852_));
 sky130_fd_sc_hd__o21ai_4 _16521_ (.A1(_01852_),
    .A2(_01728_),
    .B1(_01820_),
    .Y(_01853_));
 sky130_fd_sc_hd__inv_2 _16522_ (.A(\CPU_Xreg_value_a4[14][6] ),
    .Y(_01854_));
 sky130_fd_sc_hd__buf_2 _16523_ (.A(_01677_),
    .X(_01855_));
 sky130_fd_sc_hd__inv_2 _16524_ (.A(\CPU_Xreg_value_a4[3][6] ),
    .Y(_01856_));
 sky130_fd_sc_hd__buf_2 _16525_ (.A(_01680_),
    .X(_01857_));
 sky130_fd_sc_hd__o22a_4 _16526_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01856_),
    .B2(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__inv_2 _16527_ (.A(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__or4_4 _16528_ (.A(_01845_),
    .B(_01851_),
    .C(_01853_),
    .D(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__inv_2 _16529_ (.A(\CPU_Xreg_value_a4[1][6] ),
    .Y(_01861_));
 sky130_fd_sc_hd__buf_2 _16530_ (.A(_01685_),
    .X(_01862_));
 sky130_fd_sc_hd__inv_2 _16531_ (.A(\CPU_Xreg_value_a4[4][6] ),
    .Y(_01863_));
 sky130_fd_sc_hd__buf_2 _16532_ (.A(_01689_),
    .X(_01864_));
 sky130_fd_sc_hd__o22a_4 _16533_ (.A1(_01861_),
    .A2(_01862_),
    .B1(_01863_),
    .B2(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__inv_2 _16534_ (.A(\CPU_Xreg_value_a4[6][6] ),
    .Y(_01866_));
 sky130_fd_sc_hd__buf_2 _16535_ (.A(_01694_),
    .X(_01867_));
 sky130_fd_sc_hd__inv_2 _16536_ (.A(\CPU_Xreg_value_a4[11][6] ),
    .Y(_01868_));
 sky130_fd_sc_hd__buf_2 _16537_ (.A(_01697_),
    .X(_01869_));
 sky130_fd_sc_hd__o22a_4 _16538_ (.A1(_01866_),
    .A2(_01867_),
    .B1(_01868_),
    .B2(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__inv_2 _16539_ (.A(\CPU_Xreg_value_a4[15][6] ),
    .Y(_01871_));
 sky130_fd_sc_hd__buf_2 _16540_ (.A(_01701_),
    .X(_01872_));
 sky130_fd_sc_hd__inv_2 _16541_ (.A(\CPU_Xreg_value_a4[10][6] ),
    .Y(_01873_));
 sky130_fd_sc_hd__buf_2 _16542_ (.A(_01705_),
    .X(_01874_));
 sky130_fd_sc_hd__o22a_4 _16543_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01873_),
    .B2(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__inv_2 _16544_ (.A(\CPU_Xreg_value_a4[9][6] ),
    .Y(_01876_));
 sky130_fd_sc_hd__buf_2 _16545_ (.A(_01709_),
    .X(_01877_));
 sky130_fd_sc_hd__inv_2 _16546_ (.A(\CPU_Xreg_value_a4[7][6] ),
    .Y(_01878_));
 sky130_fd_sc_hd__buf_2 _16547_ (.A(_01712_),
    .X(_01879_));
 sky130_fd_sc_hd__o22a_4 _16548_ (.A1(_01876_),
    .A2(_01877_),
    .B1(_01878_),
    .B2(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__and4_4 _16549_ (.A(_01865_),
    .B(_01870_),
    .C(_01875_),
    .D(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__inv_2 _16550_ (.A(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__o22a_4 _16551_ (.A1(\CPU_Xreg_value_a4[0][6] ),
    .A2(_01718_),
    .B1(_01860_),
    .B2(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__o22a_4 _16552_ (.A1(_06826_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_01883_),
    .X(\CPU_src1_value_a2[6] ));
 sky130_fd_sc_hd__buf_2 _16553_ (.A(_01653_),
    .X(_01884_));
 sky130_fd_sc_hd__inv_2 _16554_ (.A(\CPU_Xreg_value_a4[8][7] ),
    .Y(_01885_));
 sky130_fd_sc_hd__buf_2 _16555_ (.A(_01657_),
    .X(_01886_));
 sky130_fd_sc_hd__buf_2 _16556_ (.A(_01721_),
    .X(_01887_));
 sky130_fd_sc_hd__a2bb2o_4 _16557_ (.A1_N(_01885_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][7] ),
    .B2(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__inv_2 _16558_ (.A(\CPU_Xreg_value_a4[5][7] ),
    .Y(_01889_));
 sky130_fd_sc_hd__inv_2 _16559_ (.A(\CPU_Xreg_value_a4[12][7] ),
    .Y(_01890_));
 sky130_fd_sc_hd__o22a_4 _16560_ (.A1(_01889_),
    .A2(_01847_),
    .B1(_01890_),
    .B2(_01849_),
    .X(_01891_));
 sky130_fd_sc_hd__inv_2 _16561_ (.A(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__inv_2 _16562_ (.A(\CPU_Xreg_value_a4[2][7] ),
    .Y(_01893_));
 sky130_fd_sc_hd__buf_2 _16563_ (.A(_01673_),
    .X(_01894_));
 sky130_fd_sc_hd__o21ai_4 _16564_ (.A1(_01893_),
    .A2(_01894_),
    .B1(_01820_),
    .Y(_01895_));
 sky130_fd_sc_hd__inv_2 _16565_ (.A(\CPU_Xreg_value_a4[14][7] ),
    .Y(_01896_));
 sky130_fd_sc_hd__inv_2 _16566_ (.A(\CPU_Xreg_value_a4[3][7] ),
    .Y(_01897_));
 sky130_fd_sc_hd__o22a_4 _16567_ (.A1(_01896_),
    .A2(_01855_),
    .B1(_01897_),
    .B2(_01857_),
    .X(_01898_));
 sky130_fd_sc_hd__inv_2 _16568_ (.A(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__or4_4 _16569_ (.A(_01888_),
    .B(_01892_),
    .C(_01895_),
    .D(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__inv_2 _16570_ (.A(\CPU_Xreg_value_a4[1][7] ),
    .Y(_01901_));
 sky130_fd_sc_hd__inv_2 _16571_ (.A(\CPU_Xreg_value_a4[4][7] ),
    .Y(_01902_));
 sky130_fd_sc_hd__o22a_4 _16572_ (.A1(_01901_),
    .A2(_01862_),
    .B1(_01902_),
    .B2(_01864_),
    .X(_01903_));
 sky130_fd_sc_hd__inv_2 _16573_ (.A(\CPU_Xreg_value_a4[6][7] ),
    .Y(_01904_));
 sky130_fd_sc_hd__inv_2 _16574_ (.A(\CPU_Xreg_value_a4[11][7] ),
    .Y(_01905_));
 sky130_fd_sc_hd__o22a_4 _16575_ (.A1(_01904_),
    .A2(_01867_),
    .B1(_01905_),
    .B2(_01869_),
    .X(_01906_));
 sky130_fd_sc_hd__inv_2 _16576_ (.A(\CPU_Xreg_value_a4[15][7] ),
    .Y(_01907_));
 sky130_fd_sc_hd__inv_2 _16577_ (.A(\CPU_Xreg_value_a4[10][7] ),
    .Y(_01908_));
 sky130_fd_sc_hd__o22a_4 _16578_ (.A1(_01907_),
    .A2(_01872_),
    .B1(_01908_),
    .B2(_01874_),
    .X(_01909_));
 sky130_fd_sc_hd__inv_2 _16579_ (.A(\CPU_Xreg_value_a4[9][7] ),
    .Y(_01910_));
 sky130_fd_sc_hd__inv_2 _16580_ (.A(\CPU_Xreg_value_a4[7][7] ),
    .Y(_01911_));
 sky130_fd_sc_hd__o22a_4 _16581_ (.A1(_01910_),
    .A2(_01877_),
    .B1(_01911_),
    .B2(_01879_),
    .X(_01912_));
 sky130_fd_sc_hd__and4_4 _16582_ (.A(_01903_),
    .B(_01906_),
    .C(_01909_),
    .D(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__inv_2 _16583_ (.A(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__o22a_4 _16584_ (.A1(\CPU_Xreg_value_a4[0][7] ),
    .A2(_01884_),
    .B1(_01900_),
    .B2(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__o22a_4 _16585_ (.A1(_06818_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_01915_),
    .X(\CPU_src1_value_a2[7] ));
 sky130_fd_sc_hd__inv_2 _16586_ (.A(\CPU_Xreg_value_a4[8][8] ),
    .Y(_01916_));
 sky130_fd_sc_hd__a2bb2o_4 _16587_ (.A1_N(_01916_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][8] ),
    .B2(_01887_),
    .X(_01917_));
 sky130_fd_sc_hd__inv_2 _16588_ (.A(\CPU_Xreg_value_a4[5][8] ),
    .Y(_01918_));
 sky130_fd_sc_hd__inv_2 _16589_ (.A(\CPU_Xreg_value_a4[12][8] ),
    .Y(_01919_));
 sky130_fd_sc_hd__o22a_4 _16590_ (.A1(_01918_),
    .A2(_01847_),
    .B1(_01919_),
    .B2(_01849_),
    .X(_01920_));
 sky130_fd_sc_hd__inv_2 _16591_ (.A(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__inv_2 _16592_ (.A(\CPU_Xreg_value_a4[2][8] ),
    .Y(_01922_));
 sky130_fd_sc_hd__o21ai_4 _16593_ (.A1(_01922_),
    .A2(_01894_),
    .B1(_01820_),
    .Y(_01923_));
 sky130_fd_sc_hd__inv_2 _16594_ (.A(\CPU_Xreg_value_a4[14][8] ),
    .Y(_01924_));
 sky130_fd_sc_hd__inv_2 _16595_ (.A(\CPU_Xreg_value_a4[3][8] ),
    .Y(_01925_));
 sky130_fd_sc_hd__o22a_4 _16596_ (.A1(_01924_),
    .A2(_01855_),
    .B1(_01925_),
    .B2(_01857_),
    .X(_01926_));
 sky130_fd_sc_hd__inv_2 _16597_ (.A(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__or4_4 _16598_ (.A(_01917_),
    .B(_01921_),
    .C(_01923_),
    .D(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__inv_2 _16599_ (.A(\CPU_Xreg_value_a4[1][8] ),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _16600_ (.A(\CPU_Xreg_value_a4[4][8] ),
    .Y(_01930_));
 sky130_fd_sc_hd__o22a_4 _16601_ (.A1(_01929_),
    .A2(_01862_),
    .B1(_01930_),
    .B2(_01864_),
    .X(_01931_));
 sky130_fd_sc_hd__inv_2 _16602_ (.A(\CPU_Xreg_value_a4[6][8] ),
    .Y(_01932_));
 sky130_fd_sc_hd__inv_2 _16603_ (.A(\CPU_Xreg_value_a4[11][8] ),
    .Y(_01933_));
 sky130_fd_sc_hd__o22a_4 _16604_ (.A1(_01932_),
    .A2(_01867_),
    .B1(_01933_),
    .B2(_01869_),
    .X(_01934_));
 sky130_fd_sc_hd__inv_2 _16605_ (.A(\CPU_Xreg_value_a4[15][8] ),
    .Y(_01935_));
 sky130_fd_sc_hd__inv_2 _16606_ (.A(\CPU_Xreg_value_a4[10][8] ),
    .Y(_01936_));
 sky130_fd_sc_hd__o22a_4 _16607_ (.A1(_01935_),
    .A2(_01872_),
    .B1(_01936_),
    .B2(_01874_),
    .X(_01937_));
 sky130_fd_sc_hd__inv_2 _16608_ (.A(\CPU_Xreg_value_a4[9][8] ),
    .Y(_01938_));
 sky130_fd_sc_hd__inv_2 _16609_ (.A(\CPU_Xreg_value_a4[7][8] ),
    .Y(_01939_));
 sky130_fd_sc_hd__o22a_4 _16610_ (.A1(_01938_),
    .A2(_01877_),
    .B1(_01939_),
    .B2(_01879_),
    .X(_01940_));
 sky130_fd_sc_hd__and4_4 _16611_ (.A(_01931_),
    .B(_01934_),
    .C(_01937_),
    .D(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__inv_2 _16612_ (.A(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__o22a_4 _16613_ (.A1(\CPU_Xreg_value_a4[0][8] ),
    .A2(_01884_),
    .B1(_01928_),
    .B2(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__o22a_4 _16614_ (.A1(_06797_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_01943_),
    .X(\CPU_src1_value_a2[8] ));
 sky130_fd_sc_hd__inv_2 _16615_ (.A(\CPU_Xreg_value_a4[8][9] ),
    .Y(_01944_));
 sky130_fd_sc_hd__a2bb2o_4 _16616_ (.A1_N(_01944_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][9] ),
    .B2(_01887_),
    .X(_01945_));
 sky130_fd_sc_hd__inv_2 _16617_ (.A(\CPU_Xreg_value_a4[5][9] ),
    .Y(_01946_));
 sky130_fd_sc_hd__inv_2 _16618_ (.A(\CPU_Xreg_value_a4[12][9] ),
    .Y(_01947_));
 sky130_fd_sc_hd__o22a_4 _16619_ (.A1(_01946_),
    .A2(_01847_),
    .B1(_01947_),
    .B2(_01849_),
    .X(_01948_));
 sky130_fd_sc_hd__inv_2 _16620_ (.A(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__inv_2 _16621_ (.A(\CPU_Xreg_value_a4[2][9] ),
    .Y(_01950_));
 sky130_fd_sc_hd__o21ai_4 _16622_ (.A1(_01950_),
    .A2(_01894_),
    .B1(_01820_),
    .Y(_01951_));
 sky130_fd_sc_hd__inv_2 _16623_ (.A(\CPU_Xreg_value_a4[14][9] ),
    .Y(_01952_));
 sky130_fd_sc_hd__inv_2 _16624_ (.A(\CPU_Xreg_value_a4[3][9] ),
    .Y(_01953_));
 sky130_fd_sc_hd__o22a_4 _16625_ (.A1(_01952_),
    .A2(_01855_),
    .B1(_01953_),
    .B2(_01857_),
    .X(_01954_));
 sky130_fd_sc_hd__inv_2 _16626_ (.A(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__or4_4 _16627_ (.A(_01945_),
    .B(_01949_),
    .C(_01951_),
    .D(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__inv_2 _16628_ (.A(\CPU_Xreg_value_a4[1][9] ),
    .Y(_01957_));
 sky130_fd_sc_hd__inv_2 _16629_ (.A(\CPU_Xreg_value_a4[4][9] ),
    .Y(_01958_));
 sky130_fd_sc_hd__o22a_4 _16630_ (.A1(_01957_),
    .A2(_01862_),
    .B1(_01958_),
    .B2(_01864_),
    .X(_01959_));
 sky130_fd_sc_hd__inv_2 _16631_ (.A(\CPU_Xreg_value_a4[6][9] ),
    .Y(_01960_));
 sky130_fd_sc_hd__inv_2 _16632_ (.A(\CPU_Xreg_value_a4[11][9] ),
    .Y(_01961_));
 sky130_fd_sc_hd__o22a_4 _16633_ (.A1(_01960_),
    .A2(_01867_),
    .B1(_01961_),
    .B2(_01869_),
    .X(_01962_));
 sky130_fd_sc_hd__inv_2 _16634_ (.A(\CPU_Xreg_value_a4[15][9] ),
    .Y(_01963_));
 sky130_fd_sc_hd__inv_2 _16635_ (.A(\CPU_Xreg_value_a4[10][9] ),
    .Y(_01964_));
 sky130_fd_sc_hd__o22a_4 _16636_ (.A1(_01963_),
    .A2(_01872_),
    .B1(_01964_),
    .B2(_01874_),
    .X(_01965_));
 sky130_fd_sc_hd__inv_2 _16637_ (.A(\CPU_Xreg_value_a4[9][9] ),
    .Y(_01966_));
 sky130_fd_sc_hd__inv_2 _16638_ (.A(\CPU_Xreg_value_a4[7][9] ),
    .Y(_01967_));
 sky130_fd_sc_hd__o22a_4 _16639_ (.A1(_01966_),
    .A2(_01877_),
    .B1(_01967_),
    .B2(_01879_),
    .X(_01968_));
 sky130_fd_sc_hd__and4_4 _16640_ (.A(_01959_),
    .B(_01962_),
    .C(_01965_),
    .D(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__inv_2 _16641_ (.A(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__o22a_4 _16642_ (.A1(\CPU_Xreg_value_a4[0][9] ),
    .A2(_01884_),
    .B1(_01956_),
    .B2(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__o22a_4 _16643_ (.A1(_06789_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_01971_),
    .X(\CPU_src1_value_a2[9] ));
 sky130_fd_sc_hd__inv_2 _16644_ (.A(\CPU_Xreg_value_a4[8][10] ),
    .Y(_01972_));
 sky130_fd_sc_hd__a2bb2o_4 _16645_ (.A1_N(_01972_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][10] ),
    .B2(_01887_),
    .X(_01973_));
 sky130_fd_sc_hd__inv_2 _16646_ (.A(\CPU_Xreg_value_a4[5][10] ),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _16647_ (.A(\CPU_Xreg_value_a4[12][10] ),
    .Y(_01975_));
 sky130_fd_sc_hd__o22a_4 _16648_ (.A1(_01974_),
    .A2(_01847_),
    .B1(_01975_),
    .B2(_01849_),
    .X(_01976_));
 sky130_fd_sc_hd__inv_2 _16649_ (.A(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__inv_2 _16650_ (.A(\CPU_Xreg_value_a4[2][10] ),
    .Y(_01978_));
 sky130_fd_sc_hd__o21ai_4 _16651_ (.A1(_01978_),
    .A2(_01894_),
    .B1(_01820_),
    .Y(_01979_));
 sky130_fd_sc_hd__inv_2 _16652_ (.A(\CPU_Xreg_value_a4[14][10] ),
    .Y(_01980_));
 sky130_fd_sc_hd__inv_2 _16653_ (.A(\CPU_Xreg_value_a4[3][10] ),
    .Y(_01981_));
 sky130_fd_sc_hd__o22a_4 _16654_ (.A1(_01980_),
    .A2(_01855_),
    .B1(_01981_),
    .B2(_01857_),
    .X(_01982_));
 sky130_fd_sc_hd__inv_2 _16655_ (.A(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__or4_4 _16656_ (.A(_01973_),
    .B(_01977_),
    .C(_01979_),
    .D(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__inv_2 _16657_ (.A(\CPU_Xreg_value_a4[1][10] ),
    .Y(_01985_));
 sky130_fd_sc_hd__inv_2 _16658_ (.A(\CPU_Xreg_value_a4[4][10] ),
    .Y(_01986_));
 sky130_fd_sc_hd__o22a_4 _16659_ (.A1(_01985_),
    .A2(_01862_),
    .B1(_01986_),
    .B2(_01864_),
    .X(_01987_));
 sky130_fd_sc_hd__inv_2 _16660_ (.A(\CPU_Xreg_value_a4[6][10] ),
    .Y(_01988_));
 sky130_fd_sc_hd__inv_2 _16661_ (.A(\CPU_Xreg_value_a4[11][10] ),
    .Y(_01989_));
 sky130_fd_sc_hd__o22a_4 _16662_ (.A1(_01988_),
    .A2(_01867_),
    .B1(_01989_),
    .B2(_01869_),
    .X(_01990_));
 sky130_fd_sc_hd__inv_2 _16663_ (.A(\CPU_Xreg_value_a4[15][10] ),
    .Y(_01991_));
 sky130_fd_sc_hd__inv_2 _16664_ (.A(\CPU_Xreg_value_a4[10][10] ),
    .Y(_01992_));
 sky130_fd_sc_hd__o22a_4 _16665_ (.A1(_01991_),
    .A2(_01872_),
    .B1(_01992_),
    .B2(_01874_),
    .X(_01993_));
 sky130_fd_sc_hd__inv_2 _16666_ (.A(\CPU_Xreg_value_a4[9][10] ),
    .Y(_01994_));
 sky130_fd_sc_hd__inv_2 _16667_ (.A(\CPU_Xreg_value_a4[7][10] ),
    .Y(_01995_));
 sky130_fd_sc_hd__o22a_4 _16668_ (.A1(_01994_),
    .A2(_01877_),
    .B1(_01995_),
    .B2(_01879_),
    .X(_01996_));
 sky130_fd_sc_hd__and4_4 _16669_ (.A(_01987_),
    .B(_01990_),
    .C(_01993_),
    .D(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__inv_2 _16670_ (.A(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o22a_4 _16671_ (.A1(\CPU_Xreg_value_a4[0][10] ),
    .A2(_01884_),
    .B1(_01984_),
    .B2(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__o22a_4 _16672_ (.A1(_06776_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_01999_),
    .X(\CPU_src1_value_a2[10] ));
 sky130_fd_sc_hd__inv_2 _16673_ (.A(\CPU_Xreg_value_a4[8][11] ),
    .Y(_02000_));
 sky130_fd_sc_hd__a2bb2o_4 _16674_ (.A1_N(_02000_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][11] ),
    .B2(_01887_),
    .X(_02001_));
 sky130_fd_sc_hd__inv_2 _16675_ (.A(\CPU_Xreg_value_a4[5][11] ),
    .Y(_02002_));
 sky130_fd_sc_hd__inv_2 _16676_ (.A(\CPU_Xreg_value_a4[12][11] ),
    .Y(_02003_));
 sky130_fd_sc_hd__o22a_4 _16677_ (.A1(_02002_),
    .A2(_01847_),
    .B1(_02003_),
    .B2(_01849_),
    .X(_02004_));
 sky130_fd_sc_hd__inv_2 _16678_ (.A(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__inv_2 _16679_ (.A(\CPU_Xreg_value_a4[2][11] ),
    .Y(_02006_));
 sky130_fd_sc_hd__buf_2 _16680_ (.A(_01650_),
    .X(_02007_));
 sky130_fd_sc_hd__o21ai_4 _16681_ (.A1(_02006_),
    .A2(_01894_),
    .B1(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__inv_2 _16682_ (.A(\CPU_Xreg_value_a4[14][11] ),
    .Y(_02009_));
 sky130_fd_sc_hd__inv_2 _16683_ (.A(\CPU_Xreg_value_a4[3][11] ),
    .Y(_02010_));
 sky130_fd_sc_hd__o22a_4 _16684_ (.A1(_02009_),
    .A2(_01855_),
    .B1(_02010_),
    .B2(_01857_),
    .X(_02011_));
 sky130_fd_sc_hd__inv_2 _16685_ (.A(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__or4_4 _16686_ (.A(_02001_),
    .B(_02005_),
    .C(_02008_),
    .D(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__inv_2 _16687_ (.A(\CPU_Xreg_value_a4[1][11] ),
    .Y(_02014_));
 sky130_fd_sc_hd__inv_2 _16688_ (.A(\CPU_Xreg_value_a4[4][11] ),
    .Y(_02015_));
 sky130_fd_sc_hd__o22a_4 _16689_ (.A1(_02014_),
    .A2(_01862_),
    .B1(_02015_),
    .B2(_01864_),
    .X(_02016_));
 sky130_fd_sc_hd__inv_2 _16690_ (.A(\CPU_Xreg_value_a4[6][11] ),
    .Y(_02017_));
 sky130_fd_sc_hd__inv_2 _16691_ (.A(\CPU_Xreg_value_a4[11][11] ),
    .Y(_02018_));
 sky130_fd_sc_hd__o22a_4 _16692_ (.A1(_02017_),
    .A2(_01867_),
    .B1(_02018_),
    .B2(_01869_),
    .X(_02019_));
 sky130_fd_sc_hd__inv_2 _16693_ (.A(\CPU_Xreg_value_a4[15][11] ),
    .Y(_02020_));
 sky130_fd_sc_hd__inv_2 _16694_ (.A(\CPU_Xreg_value_a4[10][11] ),
    .Y(_02021_));
 sky130_fd_sc_hd__o22a_4 _16695_ (.A1(_02020_),
    .A2(_01872_),
    .B1(_02021_),
    .B2(_01874_),
    .X(_02022_));
 sky130_fd_sc_hd__inv_2 _16696_ (.A(\CPU_Xreg_value_a4[9][11] ),
    .Y(_02023_));
 sky130_fd_sc_hd__inv_2 _16697_ (.A(\CPU_Xreg_value_a4[7][11] ),
    .Y(_02024_));
 sky130_fd_sc_hd__o22a_4 _16698_ (.A1(_02023_),
    .A2(_01877_),
    .B1(_02024_),
    .B2(_01879_),
    .X(_02025_));
 sky130_fd_sc_hd__and4_4 _16699_ (.A(_02016_),
    .B(_02019_),
    .C(_02022_),
    .D(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__inv_2 _16700_ (.A(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__o22a_4 _16701_ (.A1(\CPU_Xreg_value_a4[0][11] ),
    .A2(_01884_),
    .B1(_02013_),
    .B2(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__o22a_4 _16702_ (.A1(_06768_),
    .A2(_01842_),
    .B1(_01843_),
    .B2(_02028_),
    .X(\CPU_src1_value_a2[11] ));
 sky130_fd_sc_hd__buf_2 _16703_ (.A(_01644_),
    .X(_02029_));
 sky130_fd_sc_hd__buf_2 _16704_ (.A(_01647_),
    .X(_02030_));
 sky130_fd_sc_hd__inv_2 _16705_ (.A(\CPU_Xreg_value_a4[8][12] ),
    .Y(_02031_));
 sky130_fd_sc_hd__a2bb2o_4 _16706_ (.A1_N(_02031_),
    .A2_N(_01886_),
    .B1(\CPU_Xreg_value_a4[13][12] ),
    .B2(_01887_),
    .X(_02032_));
 sky130_fd_sc_hd__inv_2 _16707_ (.A(\CPU_Xreg_value_a4[5][12] ),
    .Y(_02033_));
 sky130_fd_sc_hd__buf_2 _16708_ (.A(_01664_),
    .X(_02034_));
 sky130_fd_sc_hd__inv_2 _16709_ (.A(\CPU_Xreg_value_a4[12][12] ),
    .Y(_02035_));
 sky130_fd_sc_hd__buf_2 _16710_ (.A(_01668_),
    .X(_02036_));
 sky130_fd_sc_hd__o22a_4 _16711_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_02035_),
    .B2(_02036_),
    .X(_02037_));
 sky130_fd_sc_hd__inv_2 _16712_ (.A(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__inv_2 _16713_ (.A(\CPU_Xreg_value_a4[2][12] ),
    .Y(_02039_));
 sky130_fd_sc_hd__o21ai_4 _16714_ (.A1(_02039_),
    .A2(_01894_),
    .B1(_02007_),
    .Y(_02040_));
 sky130_fd_sc_hd__inv_2 _16715_ (.A(\CPU_Xreg_value_a4[14][12] ),
    .Y(_02041_));
 sky130_fd_sc_hd__buf_2 _16716_ (.A(_01677_),
    .X(_02042_));
 sky130_fd_sc_hd__inv_2 _16717_ (.A(\CPU_Xreg_value_a4[3][12] ),
    .Y(_02043_));
 sky130_fd_sc_hd__buf_2 _16718_ (.A(_01680_),
    .X(_02044_));
 sky130_fd_sc_hd__o22a_4 _16719_ (.A1(_02041_),
    .A2(_02042_),
    .B1(_02043_),
    .B2(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__inv_2 _16720_ (.A(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__or4_4 _16721_ (.A(_02032_),
    .B(_02038_),
    .C(_02040_),
    .D(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__inv_2 _16722_ (.A(\CPU_Xreg_value_a4[1][12] ),
    .Y(_02048_));
 sky130_fd_sc_hd__buf_2 _16723_ (.A(_01685_),
    .X(_02049_));
 sky130_fd_sc_hd__inv_2 _16724_ (.A(\CPU_Xreg_value_a4[4][12] ),
    .Y(_02050_));
 sky130_fd_sc_hd__buf_2 _16725_ (.A(_01689_),
    .X(_02051_));
 sky130_fd_sc_hd__o22a_4 _16726_ (.A1(_02048_),
    .A2(_02049_),
    .B1(_02050_),
    .B2(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__inv_2 _16727_ (.A(\CPU_Xreg_value_a4[6][12] ),
    .Y(_02053_));
 sky130_fd_sc_hd__buf_2 _16728_ (.A(_01694_),
    .X(_02054_));
 sky130_fd_sc_hd__inv_2 _16729_ (.A(\CPU_Xreg_value_a4[11][12] ),
    .Y(_02055_));
 sky130_fd_sc_hd__buf_2 _16730_ (.A(_01697_),
    .X(_02056_));
 sky130_fd_sc_hd__o22a_4 _16731_ (.A1(_02053_),
    .A2(_02054_),
    .B1(_02055_),
    .B2(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__inv_2 _16732_ (.A(\CPU_Xreg_value_a4[15][12] ),
    .Y(_02058_));
 sky130_fd_sc_hd__buf_2 _16733_ (.A(_01701_),
    .X(_02059_));
 sky130_fd_sc_hd__inv_2 _16734_ (.A(\CPU_Xreg_value_a4[10][12] ),
    .Y(_02060_));
 sky130_fd_sc_hd__buf_2 _16735_ (.A(_01705_),
    .X(_02061_));
 sky130_fd_sc_hd__o22a_4 _16736_ (.A1(_02058_),
    .A2(_02059_),
    .B1(_02060_),
    .B2(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__inv_2 _16737_ (.A(\CPU_Xreg_value_a4[9][12] ),
    .Y(_02063_));
 sky130_fd_sc_hd__buf_2 _16738_ (.A(_01709_),
    .X(_02064_));
 sky130_fd_sc_hd__inv_2 _16739_ (.A(\CPU_Xreg_value_a4[7][12] ),
    .Y(_02065_));
 sky130_fd_sc_hd__buf_2 _16740_ (.A(_01712_),
    .X(_02066_));
 sky130_fd_sc_hd__o22a_4 _16741_ (.A1(_02063_),
    .A2(_02064_),
    .B1(_02065_),
    .B2(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__and4_4 _16742_ (.A(_02052_),
    .B(_02057_),
    .C(_02062_),
    .D(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__inv_2 _16743_ (.A(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__o22a_4 _16744_ (.A1(\CPU_Xreg_value_a4[0][12] ),
    .A2(_01884_),
    .B1(_02047_),
    .B2(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__o22a_4 _16745_ (.A1(_06750_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02070_),
    .X(\CPU_src1_value_a2[12] ));
 sky130_fd_sc_hd__buf_2 _16746_ (.A(_01653_),
    .X(_02071_));
 sky130_fd_sc_hd__inv_2 _16747_ (.A(\CPU_Xreg_value_a4[8][13] ),
    .Y(_02072_));
 sky130_fd_sc_hd__buf_2 _16748_ (.A(_01657_),
    .X(_02073_));
 sky130_fd_sc_hd__buf_2 _16749_ (.A(_01721_),
    .X(_02074_));
 sky130_fd_sc_hd__a2bb2o_4 _16750_ (.A1_N(_02072_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][13] ),
    .B2(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__inv_2 _16751_ (.A(\CPU_Xreg_value_a4[5][13] ),
    .Y(_02076_));
 sky130_fd_sc_hd__inv_2 _16752_ (.A(\CPU_Xreg_value_a4[12][13] ),
    .Y(_02077_));
 sky130_fd_sc_hd__o22a_4 _16753_ (.A1(_02076_),
    .A2(_02034_),
    .B1(_02077_),
    .B2(_02036_),
    .X(_02078_));
 sky130_fd_sc_hd__inv_2 _16754_ (.A(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__inv_2 _16755_ (.A(\CPU_Xreg_value_a4[2][13] ),
    .Y(_02080_));
 sky130_fd_sc_hd__buf_2 _16756_ (.A(_01673_),
    .X(_02081_));
 sky130_fd_sc_hd__o21ai_4 _16757_ (.A1(_02080_),
    .A2(_02081_),
    .B1(_02007_),
    .Y(_02082_));
 sky130_fd_sc_hd__inv_2 _16758_ (.A(\CPU_Xreg_value_a4[14][13] ),
    .Y(_02083_));
 sky130_fd_sc_hd__inv_2 _16759_ (.A(\CPU_Xreg_value_a4[3][13] ),
    .Y(_02084_));
 sky130_fd_sc_hd__o22a_4 _16760_ (.A1(_02083_),
    .A2(_02042_),
    .B1(_02084_),
    .B2(_02044_),
    .X(_02085_));
 sky130_fd_sc_hd__inv_2 _16761_ (.A(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__or4_4 _16762_ (.A(_02075_),
    .B(_02079_),
    .C(_02082_),
    .D(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__inv_2 _16763_ (.A(\CPU_Xreg_value_a4[1][13] ),
    .Y(_02088_));
 sky130_fd_sc_hd__inv_2 _16764_ (.A(\CPU_Xreg_value_a4[4][13] ),
    .Y(_02089_));
 sky130_fd_sc_hd__o22a_4 _16765_ (.A1(_02088_),
    .A2(_02049_),
    .B1(_02089_),
    .B2(_02051_),
    .X(_02090_));
 sky130_fd_sc_hd__inv_2 _16766_ (.A(\CPU_Xreg_value_a4[6][13] ),
    .Y(_02091_));
 sky130_fd_sc_hd__inv_2 _16767_ (.A(\CPU_Xreg_value_a4[11][13] ),
    .Y(_02092_));
 sky130_fd_sc_hd__o22a_4 _16768_ (.A1(_02091_),
    .A2(_02054_),
    .B1(_02092_),
    .B2(_02056_),
    .X(_02093_));
 sky130_fd_sc_hd__inv_2 _16769_ (.A(\CPU_Xreg_value_a4[15][13] ),
    .Y(_02094_));
 sky130_fd_sc_hd__inv_2 _16770_ (.A(\CPU_Xreg_value_a4[10][13] ),
    .Y(_02095_));
 sky130_fd_sc_hd__o22a_4 _16771_ (.A1(_02094_),
    .A2(_02059_),
    .B1(_02095_),
    .B2(_02061_),
    .X(_02096_));
 sky130_fd_sc_hd__inv_2 _16772_ (.A(\CPU_Xreg_value_a4[9][13] ),
    .Y(_02097_));
 sky130_fd_sc_hd__inv_2 _16773_ (.A(\CPU_Xreg_value_a4[7][13] ),
    .Y(_02098_));
 sky130_fd_sc_hd__o22a_4 _16774_ (.A1(_02097_),
    .A2(_02064_),
    .B1(_02098_),
    .B2(_02066_),
    .X(_02099_));
 sky130_fd_sc_hd__and4_4 _16775_ (.A(_02090_),
    .B(_02093_),
    .C(_02096_),
    .D(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__inv_2 _16776_ (.A(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__o22a_4 _16777_ (.A1(\CPU_Xreg_value_a4[0][13] ),
    .A2(_02071_),
    .B1(_02087_),
    .B2(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__o22a_4 _16778_ (.A1(_06741_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02102_),
    .X(\CPU_src1_value_a2[13] ));
 sky130_fd_sc_hd__inv_2 _16779_ (.A(\CPU_Xreg_value_a4[8][14] ),
    .Y(_02103_));
 sky130_fd_sc_hd__a2bb2o_4 _16780_ (.A1_N(_02103_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][14] ),
    .B2(_02074_),
    .X(_02104_));
 sky130_fd_sc_hd__inv_2 _16781_ (.A(\CPU_Xreg_value_a4[5][14] ),
    .Y(_02105_));
 sky130_fd_sc_hd__inv_2 _16782_ (.A(\CPU_Xreg_value_a4[12][14] ),
    .Y(_02106_));
 sky130_fd_sc_hd__o22a_4 _16783_ (.A1(_02105_),
    .A2(_02034_),
    .B1(_02106_),
    .B2(_02036_),
    .X(_02107_));
 sky130_fd_sc_hd__inv_2 _16784_ (.A(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__inv_2 _16785_ (.A(\CPU_Xreg_value_a4[2][14] ),
    .Y(_02109_));
 sky130_fd_sc_hd__o21ai_4 _16786_ (.A1(_02109_),
    .A2(_02081_),
    .B1(_02007_),
    .Y(_02110_));
 sky130_fd_sc_hd__inv_2 _16787_ (.A(\CPU_Xreg_value_a4[14][14] ),
    .Y(_02111_));
 sky130_fd_sc_hd__inv_2 _16788_ (.A(\CPU_Xreg_value_a4[3][14] ),
    .Y(_02112_));
 sky130_fd_sc_hd__o22a_4 _16789_ (.A1(_02111_),
    .A2(_02042_),
    .B1(_02112_),
    .B2(_02044_),
    .X(_02113_));
 sky130_fd_sc_hd__inv_2 _16790_ (.A(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__or4_4 _16791_ (.A(_02104_),
    .B(_02108_),
    .C(_02110_),
    .D(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__inv_2 _16792_ (.A(\CPU_Xreg_value_a4[1][14] ),
    .Y(_02116_));
 sky130_fd_sc_hd__inv_2 _16793_ (.A(\CPU_Xreg_value_a4[4][14] ),
    .Y(_02117_));
 sky130_fd_sc_hd__o22a_4 _16794_ (.A1(_02116_),
    .A2(_02049_),
    .B1(_02117_),
    .B2(_02051_),
    .X(_02118_));
 sky130_fd_sc_hd__inv_2 _16795_ (.A(\CPU_Xreg_value_a4[6][14] ),
    .Y(_02119_));
 sky130_fd_sc_hd__inv_2 _16796_ (.A(\CPU_Xreg_value_a4[11][14] ),
    .Y(_02120_));
 sky130_fd_sc_hd__o22a_4 _16797_ (.A1(_02119_),
    .A2(_02054_),
    .B1(_02120_),
    .B2(_02056_),
    .X(_02121_));
 sky130_fd_sc_hd__inv_2 _16798_ (.A(\CPU_Xreg_value_a4[15][14] ),
    .Y(_02122_));
 sky130_fd_sc_hd__inv_2 _16799_ (.A(\CPU_Xreg_value_a4[10][14] ),
    .Y(_02123_));
 sky130_fd_sc_hd__o22a_4 _16800_ (.A1(_02122_),
    .A2(_02059_),
    .B1(_02123_),
    .B2(_02061_),
    .X(_02124_));
 sky130_fd_sc_hd__inv_2 _16801_ (.A(\CPU_Xreg_value_a4[9][14] ),
    .Y(_02125_));
 sky130_fd_sc_hd__inv_2 _16802_ (.A(\CPU_Xreg_value_a4[7][14] ),
    .Y(_02126_));
 sky130_fd_sc_hd__o22a_4 _16803_ (.A1(_02125_),
    .A2(_02064_),
    .B1(_02126_),
    .B2(_02066_),
    .X(_02127_));
 sky130_fd_sc_hd__and4_4 _16804_ (.A(_02118_),
    .B(_02121_),
    .C(_02124_),
    .D(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__inv_2 _16805_ (.A(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__o22a_4 _16806_ (.A1(\CPU_Xreg_value_a4[0][14] ),
    .A2(_02071_),
    .B1(_02115_),
    .B2(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__o22a_4 _16807_ (.A1(_06731_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02130_),
    .X(\CPU_src1_value_a2[14] ));
 sky130_fd_sc_hd__inv_2 _16808_ (.A(\CPU_Xreg_value_a4[8][15] ),
    .Y(_02131_));
 sky130_fd_sc_hd__a2bb2o_4 _16809_ (.A1_N(_02131_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][15] ),
    .B2(_02074_),
    .X(_02132_));
 sky130_fd_sc_hd__inv_2 _16810_ (.A(\CPU_Xreg_value_a4[5][15] ),
    .Y(_02133_));
 sky130_fd_sc_hd__inv_2 _16811_ (.A(\CPU_Xreg_value_a4[12][15] ),
    .Y(_02134_));
 sky130_fd_sc_hd__o22a_4 _16812_ (.A1(_02133_),
    .A2(_02034_),
    .B1(_02134_),
    .B2(_02036_),
    .X(_02135_));
 sky130_fd_sc_hd__inv_2 _16813_ (.A(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__inv_2 _16814_ (.A(\CPU_Xreg_value_a4[2][15] ),
    .Y(_02137_));
 sky130_fd_sc_hd__o21ai_4 _16815_ (.A1(_02137_),
    .A2(_02081_),
    .B1(_02007_),
    .Y(_02138_));
 sky130_fd_sc_hd__inv_2 _16816_ (.A(\CPU_Xreg_value_a4[14][15] ),
    .Y(_02139_));
 sky130_fd_sc_hd__inv_2 _16817_ (.A(\CPU_Xreg_value_a4[3][15] ),
    .Y(_02140_));
 sky130_fd_sc_hd__o22a_4 _16818_ (.A1(_02139_),
    .A2(_02042_),
    .B1(_02140_),
    .B2(_02044_),
    .X(_02141_));
 sky130_fd_sc_hd__inv_2 _16819_ (.A(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__or4_4 _16820_ (.A(_02132_),
    .B(_02136_),
    .C(_02138_),
    .D(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__inv_2 _16821_ (.A(\CPU_Xreg_value_a4[1][15] ),
    .Y(_02144_));
 sky130_fd_sc_hd__inv_2 _16822_ (.A(\CPU_Xreg_value_a4[4][15] ),
    .Y(_02145_));
 sky130_fd_sc_hd__o22a_4 _16823_ (.A1(_02144_),
    .A2(_02049_),
    .B1(_02145_),
    .B2(_02051_),
    .X(_02146_));
 sky130_fd_sc_hd__inv_2 _16824_ (.A(\CPU_Xreg_value_a4[6][15] ),
    .Y(_02147_));
 sky130_fd_sc_hd__inv_2 _16825_ (.A(\CPU_Xreg_value_a4[11][15] ),
    .Y(_02148_));
 sky130_fd_sc_hd__o22a_4 _16826_ (.A1(_02147_),
    .A2(_02054_),
    .B1(_02148_),
    .B2(_02056_),
    .X(_02149_));
 sky130_fd_sc_hd__inv_2 _16827_ (.A(\CPU_Xreg_value_a4[15][15] ),
    .Y(_02150_));
 sky130_fd_sc_hd__inv_2 _16828_ (.A(\CPU_Xreg_value_a4[10][15] ),
    .Y(_02151_));
 sky130_fd_sc_hd__o22a_4 _16829_ (.A1(_02150_),
    .A2(_02059_),
    .B1(_02151_),
    .B2(_02061_),
    .X(_02152_));
 sky130_fd_sc_hd__inv_2 _16830_ (.A(\CPU_Xreg_value_a4[9][15] ),
    .Y(_02153_));
 sky130_fd_sc_hd__inv_2 _16831_ (.A(\CPU_Xreg_value_a4[7][15] ),
    .Y(_02154_));
 sky130_fd_sc_hd__o22a_4 _16832_ (.A1(_02153_),
    .A2(_02064_),
    .B1(_02154_),
    .B2(_02066_),
    .X(_02155_));
 sky130_fd_sc_hd__and4_4 _16833_ (.A(_02146_),
    .B(_02149_),
    .C(_02152_),
    .D(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__inv_2 _16834_ (.A(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__o22a_4 _16835_ (.A1(\CPU_Xreg_value_a4[0][15] ),
    .A2(_02071_),
    .B1(_02143_),
    .B2(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__o22a_4 _16836_ (.A1(_06722_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02158_),
    .X(\CPU_src1_value_a2[15] ));
 sky130_fd_sc_hd__inv_2 _16837_ (.A(\CPU_Xreg_value_a4[8][16] ),
    .Y(_02159_));
 sky130_fd_sc_hd__a2bb2o_4 _16838_ (.A1_N(_02159_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][16] ),
    .B2(_02074_),
    .X(_02160_));
 sky130_fd_sc_hd__inv_2 _16839_ (.A(\CPU_Xreg_value_a4[5][16] ),
    .Y(_02161_));
 sky130_fd_sc_hd__inv_2 _16840_ (.A(\CPU_Xreg_value_a4[12][16] ),
    .Y(_02162_));
 sky130_fd_sc_hd__o22a_4 _16841_ (.A1(_02161_),
    .A2(_02034_),
    .B1(_02162_),
    .B2(_02036_),
    .X(_02163_));
 sky130_fd_sc_hd__inv_2 _16842_ (.A(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__inv_2 _16843_ (.A(\CPU_Xreg_value_a4[2][16] ),
    .Y(_02165_));
 sky130_fd_sc_hd__o21ai_4 _16844_ (.A1(_02165_),
    .A2(_02081_),
    .B1(_02007_),
    .Y(_02166_));
 sky130_fd_sc_hd__inv_2 _16845_ (.A(\CPU_Xreg_value_a4[14][16] ),
    .Y(_02167_));
 sky130_fd_sc_hd__inv_2 _16846_ (.A(\CPU_Xreg_value_a4[3][16] ),
    .Y(_02168_));
 sky130_fd_sc_hd__o22a_4 _16847_ (.A1(_02167_),
    .A2(_02042_),
    .B1(_02168_),
    .B2(_02044_),
    .X(_02169_));
 sky130_fd_sc_hd__inv_2 _16848_ (.A(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__or4_4 _16849_ (.A(_02160_),
    .B(_02164_),
    .C(_02166_),
    .D(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__inv_2 _16850_ (.A(\CPU_Xreg_value_a4[1][16] ),
    .Y(_02172_));
 sky130_fd_sc_hd__inv_2 _16851_ (.A(\CPU_Xreg_value_a4[4][16] ),
    .Y(_02173_));
 sky130_fd_sc_hd__o22a_4 _16852_ (.A1(_02172_),
    .A2(_02049_),
    .B1(_02173_),
    .B2(_02051_),
    .X(_02174_));
 sky130_fd_sc_hd__inv_2 _16853_ (.A(\CPU_Xreg_value_a4[6][16] ),
    .Y(_02175_));
 sky130_fd_sc_hd__inv_2 _16854_ (.A(\CPU_Xreg_value_a4[11][16] ),
    .Y(_02176_));
 sky130_fd_sc_hd__o22a_4 _16855_ (.A1(_02175_),
    .A2(_02054_),
    .B1(_02176_),
    .B2(_02056_),
    .X(_02177_));
 sky130_fd_sc_hd__inv_2 _16856_ (.A(\CPU_Xreg_value_a4[15][16] ),
    .Y(_02178_));
 sky130_fd_sc_hd__inv_2 _16857_ (.A(\CPU_Xreg_value_a4[10][16] ),
    .Y(_02179_));
 sky130_fd_sc_hd__o22a_4 _16858_ (.A1(_02178_),
    .A2(_02059_),
    .B1(_02179_),
    .B2(_02061_),
    .X(_02180_));
 sky130_fd_sc_hd__inv_2 _16859_ (.A(\CPU_Xreg_value_a4[9][16] ),
    .Y(_02181_));
 sky130_fd_sc_hd__inv_2 _16860_ (.A(\CPU_Xreg_value_a4[7][16] ),
    .Y(_02182_));
 sky130_fd_sc_hd__o22a_4 _16861_ (.A1(_02181_),
    .A2(_02064_),
    .B1(_02182_),
    .B2(_02066_),
    .X(_02183_));
 sky130_fd_sc_hd__and4_4 _16862_ (.A(_02174_),
    .B(_02177_),
    .C(_02180_),
    .D(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__inv_2 _16863_ (.A(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__o22a_4 _16864_ (.A1(\CPU_Xreg_value_a4[0][16] ),
    .A2(_02071_),
    .B1(_02171_),
    .B2(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__o22a_4 _16865_ (.A1(_06699_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02186_),
    .X(\CPU_src1_value_a2[16] ));
 sky130_fd_sc_hd__inv_2 _16866_ (.A(\CPU_Xreg_value_a4[8][17] ),
    .Y(_02187_));
 sky130_fd_sc_hd__a2bb2o_4 _16867_ (.A1_N(_02187_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][17] ),
    .B2(_02074_),
    .X(_02188_));
 sky130_fd_sc_hd__inv_2 _16868_ (.A(\CPU_Xreg_value_a4[5][17] ),
    .Y(_02189_));
 sky130_fd_sc_hd__inv_2 _16869_ (.A(\CPU_Xreg_value_a4[12][17] ),
    .Y(_02190_));
 sky130_fd_sc_hd__o22a_4 _16870_ (.A1(_02189_),
    .A2(_02034_),
    .B1(_02190_),
    .B2(_02036_),
    .X(_02191_));
 sky130_fd_sc_hd__inv_2 _16871_ (.A(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__inv_2 _16872_ (.A(\CPU_Xreg_value_a4[2][17] ),
    .Y(_02193_));
 sky130_fd_sc_hd__buf_2 _16873_ (.A(_01650_),
    .X(_02194_));
 sky130_fd_sc_hd__o21ai_4 _16874_ (.A1(_02193_),
    .A2(_02081_),
    .B1(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__inv_2 _16875_ (.A(\CPU_Xreg_value_a4[14][17] ),
    .Y(_02196_));
 sky130_fd_sc_hd__inv_2 _16876_ (.A(\CPU_Xreg_value_a4[3][17] ),
    .Y(_02197_));
 sky130_fd_sc_hd__o22a_4 _16877_ (.A1(_02196_),
    .A2(_02042_),
    .B1(_02197_),
    .B2(_02044_),
    .X(_02198_));
 sky130_fd_sc_hd__inv_2 _16878_ (.A(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__or4_4 _16879_ (.A(_02188_),
    .B(_02192_),
    .C(_02195_),
    .D(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__inv_2 _16880_ (.A(\CPU_Xreg_value_a4[1][17] ),
    .Y(_02201_));
 sky130_fd_sc_hd__inv_2 _16881_ (.A(\CPU_Xreg_value_a4[4][17] ),
    .Y(_02202_));
 sky130_fd_sc_hd__o22a_4 _16882_ (.A1(_02201_),
    .A2(_02049_),
    .B1(_02202_),
    .B2(_02051_),
    .X(_02203_));
 sky130_fd_sc_hd__inv_2 _16883_ (.A(\CPU_Xreg_value_a4[6][17] ),
    .Y(_02204_));
 sky130_fd_sc_hd__inv_2 _16884_ (.A(\CPU_Xreg_value_a4[11][17] ),
    .Y(_02205_));
 sky130_fd_sc_hd__o22a_4 _16885_ (.A1(_02204_),
    .A2(_02054_),
    .B1(_02205_),
    .B2(_02056_),
    .X(_02206_));
 sky130_fd_sc_hd__inv_2 _16886_ (.A(\CPU_Xreg_value_a4[15][17] ),
    .Y(_02207_));
 sky130_fd_sc_hd__inv_2 _16887_ (.A(\CPU_Xreg_value_a4[10][17] ),
    .Y(_02208_));
 sky130_fd_sc_hd__o22a_4 _16888_ (.A1(_02207_),
    .A2(_02059_),
    .B1(_02208_),
    .B2(_02061_),
    .X(_02209_));
 sky130_fd_sc_hd__inv_2 _16889_ (.A(\CPU_Xreg_value_a4[9][17] ),
    .Y(_02210_));
 sky130_fd_sc_hd__inv_2 _16890_ (.A(\CPU_Xreg_value_a4[7][17] ),
    .Y(_02211_));
 sky130_fd_sc_hd__o22a_4 _16891_ (.A1(_02210_),
    .A2(_02064_),
    .B1(_02211_),
    .B2(_02066_),
    .X(_02212_));
 sky130_fd_sc_hd__and4_4 _16892_ (.A(_02203_),
    .B(_02206_),
    .C(_02209_),
    .D(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__inv_2 _16893_ (.A(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__o22a_4 _16894_ (.A1(\CPU_Xreg_value_a4[0][17] ),
    .A2(_02071_),
    .B1(_02200_),
    .B2(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__o22a_4 _16895_ (.A1(_06690_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02215_),
    .X(\CPU_src1_value_a2[17] ));
 sky130_fd_sc_hd__buf_2 _16896_ (.A(_01644_),
    .X(_02216_));
 sky130_fd_sc_hd__buf_2 _16897_ (.A(_01647_),
    .X(_02217_));
 sky130_fd_sc_hd__inv_2 _16898_ (.A(\CPU_Xreg_value_a4[8][18] ),
    .Y(_02218_));
 sky130_fd_sc_hd__a2bb2o_4 _16899_ (.A1_N(_02218_),
    .A2_N(_02073_),
    .B1(\CPU_Xreg_value_a4[13][18] ),
    .B2(_02074_),
    .X(_02219_));
 sky130_fd_sc_hd__inv_2 _16900_ (.A(\CPU_Xreg_value_a4[5][18] ),
    .Y(_02220_));
 sky130_fd_sc_hd__buf_2 _16901_ (.A(_01664_),
    .X(_02221_));
 sky130_fd_sc_hd__inv_2 _16902_ (.A(\CPU_Xreg_value_a4[12][18] ),
    .Y(_02222_));
 sky130_fd_sc_hd__buf_2 _16903_ (.A(_01668_),
    .X(_02223_));
 sky130_fd_sc_hd__o22a_4 _16904_ (.A1(_02220_),
    .A2(_02221_),
    .B1(_02222_),
    .B2(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__inv_2 _16905_ (.A(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__inv_2 _16906_ (.A(\CPU_Xreg_value_a4[2][18] ),
    .Y(_02226_));
 sky130_fd_sc_hd__o21ai_4 _16907_ (.A1(_02226_),
    .A2(_02081_),
    .B1(_02194_),
    .Y(_02227_));
 sky130_fd_sc_hd__inv_2 _16908_ (.A(\CPU_Xreg_value_a4[14][18] ),
    .Y(_02228_));
 sky130_fd_sc_hd__buf_2 _16909_ (.A(_01677_),
    .X(_02229_));
 sky130_fd_sc_hd__inv_2 _16910_ (.A(\CPU_Xreg_value_a4[3][18] ),
    .Y(_02230_));
 sky130_fd_sc_hd__buf_2 _16911_ (.A(_01680_),
    .X(_02231_));
 sky130_fd_sc_hd__o22a_4 _16912_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02230_),
    .B2(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__inv_2 _16913_ (.A(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__or4_4 _16914_ (.A(_02219_),
    .B(_02225_),
    .C(_02227_),
    .D(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__inv_2 _16915_ (.A(\CPU_Xreg_value_a4[1][18] ),
    .Y(_02235_));
 sky130_fd_sc_hd__buf_2 _16916_ (.A(_01685_),
    .X(_02236_));
 sky130_fd_sc_hd__inv_2 _16917_ (.A(\CPU_Xreg_value_a4[4][18] ),
    .Y(_02237_));
 sky130_fd_sc_hd__buf_2 _16918_ (.A(_01689_),
    .X(_02238_));
 sky130_fd_sc_hd__o22a_4 _16919_ (.A1(_02235_),
    .A2(_02236_),
    .B1(_02237_),
    .B2(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__inv_2 _16920_ (.A(\CPU_Xreg_value_a4[6][18] ),
    .Y(_02240_));
 sky130_fd_sc_hd__buf_2 _16921_ (.A(_01694_),
    .X(_02241_));
 sky130_fd_sc_hd__inv_2 _16922_ (.A(\CPU_Xreg_value_a4[11][18] ),
    .Y(_02242_));
 sky130_fd_sc_hd__buf_2 _16923_ (.A(_01697_),
    .X(_02243_));
 sky130_fd_sc_hd__o22a_4 _16924_ (.A1(_02240_),
    .A2(_02241_),
    .B1(_02242_),
    .B2(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__inv_2 _16925_ (.A(\CPU_Xreg_value_a4[15][18] ),
    .Y(_02245_));
 sky130_fd_sc_hd__buf_2 _16926_ (.A(_01701_),
    .X(_02246_));
 sky130_fd_sc_hd__inv_2 _16927_ (.A(\CPU_Xreg_value_a4[10][18] ),
    .Y(_02247_));
 sky130_fd_sc_hd__buf_2 _16928_ (.A(_01705_),
    .X(_02248_));
 sky130_fd_sc_hd__o22a_4 _16929_ (.A1(_02245_),
    .A2(_02246_),
    .B1(_02247_),
    .B2(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__inv_2 _16930_ (.A(\CPU_Xreg_value_a4[9][18] ),
    .Y(_02250_));
 sky130_fd_sc_hd__buf_2 _16931_ (.A(_01709_),
    .X(_02251_));
 sky130_fd_sc_hd__inv_2 _16932_ (.A(\CPU_Xreg_value_a4[7][18] ),
    .Y(_02252_));
 sky130_fd_sc_hd__buf_2 _16933_ (.A(_01712_),
    .X(_02253_));
 sky130_fd_sc_hd__o22a_4 _16934_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_02252_),
    .B2(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__and4_4 _16935_ (.A(_02239_),
    .B(_02244_),
    .C(_02249_),
    .D(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__inv_2 _16936_ (.A(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__o22a_4 _16937_ (.A1(\CPU_Xreg_value_a4[0][18] ),
    .A2(_02071_),
    .B1(_02234_),
    .B2(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__o22a_4 _16938_ (.A1(_06680_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02257_),
    .X(\CPU_src1_value_a2[18] ));
 sky130_fd_sc_hd__buf_2 _16939_ (.A(_01653_),
    .X(_02258_));
 sky130_fd_sc_hd__inv_2 _16940_ (.A(\CPU_Xreg_value_a4[8][19] ),
    .Y(_02259_));
 sky130_fd_sc_hd__buf_2 _16941_ (.A(_01657_),
    .X(_02260_));
 sky130_fd_sc_hd__buf_2 _16942_ (.A(_01721_),
    .X(_02261_));
 sky130_fd_sc_hd__a2bb2o_4 _16943_ (.A1_N(_02259_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][19] ),
    .B2(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__inv_2 _16944_ (.A(\CPU_Xreg_value_a4[5][19] ),
    .Y(_02263_));
 sky130_fd_sc_hd__inv_2 _16945_ (.A(\CPU_Xreg_value_a4[12][19] ),
    .Y(_02264_));
 sky130_fd_sc_hd__o22a_4 _16946_ (.A1(_02263_),
    .A2(_02221_),
    .B1(_02264_),
    .B2(_02223_),
    .X(_02265_));
 sky130_fd_sc_hd__inv_2 _16947_ (.A(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__inv_2 _16948_ (.A(\CPU_Xreg_value_a4[2][19] ),
    .Y(_02267_));
 sky130_fd_sc_hd__buf_2 _16949_ (.A(_01673_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_4 _16950_ (.A1(_02267_),
    .A2(_02268_),
    .B1(_02194_),
    .Y(_02269_));
 sky130_fd_sc_hd__inv_2 _16951_ (.A(\CPU_Xreg_value_a4[14][19] ),
    .Y(_02270_));
 sky130_fd_sc_hd__inv_2 _16952_ (.A(\CPU_Xreg_value_a4[3][19] ),
    .Y(_02271_));
 sky130_fd_sc_hd__o22a_4 _16953_ (.A1(_02270_),
    .A2(_02229_),
    .B1(_02271_),
    .B2(_02231_),
    .X(_02272_));
 sky130_fd_sc_hd__inv_2 _16954_ (.A(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__or4_4 _16955_ (.A(_02262_),
    .B(_02266_),
    .C(_02269_),
    .D(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__inv_2 _16956_ (.A(\CPU_Xreg_value_a4[1][19] ),
    .Y(_02275_));
 sky130_fd_sc_hd__inv_2 _16957_ (.A(\CPU_Xreg_value_a4[4][19] ),
    .Y(_02276_));
 sky130_fd_sc_hd__o22a_4 _16958_ (.A1(_02275_),
    .A2(_02236_),
    .B1(_02276_),
    .B2(_02238_),
    .X(_02277_));
 sky130_fd_sc_hd__inv_2 _16959_ (.A(\CPU_Xreg_value_a4[6][19] ),
    .Y(_02278_));
 sky130_fd_sc_hd__inv_2 _16960_ (.A(\CPU_Xreg_value_a4[11][19] ),
    .Y(_02279_));
 sky130_fd_sc_hd__o22a_4 _16961_ (.A1(_02278_),
    .A2(_02241_),
    .B1(_02279_),
    .B2(_02243_),
    .X(_02280_));
 sky130_fd_sc_hd__inv_2 _16962_ (.A(\CPU_Xreg_value_a4[15][19] ),
    .Y(_02281_));
 sky130_fd_sc_hd__inv_2 _16963_ (.A(\CPU_Xreg_value_a4[10][19] ),
    .Y(_02282_));
 sky130_fd_sc_hd__o22a_4 _16964_ (.A1(_02281_),
    .A2(_02246_),
    .B1(_02282_),
    .B2(_02248_),
    .X(_02283_));
 sky130_fd_sc_hd__inv_2 _16965_ (.A(\CPU_Xreg_value_a4[9][19] ),
    .Y(_02284_));
 sky130_fd_sc_hd__inv_2 _16966_ (.A(\CPU_Xreg_value_a4[7][19] ),
    .Y(_02285_));
 sky130_fd_sc_hd__o22a_4 _16967_ (.A1(_02284_),
    .A2(_02251_),
    .B1(_02285_),
    .B2(_02253_),
    .X(_02286_));
 sky130_fd_sc_hd__and4_4 _16968_ (.A(_02277_),
    .B(_02280_),
    .C(_02283_),
    .D(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__inv_2 _16969_ (.A(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__o22a_4 _16970_ (.A1(\CPU_Xreg_value_a4[0][19] ),
    .A2(_02258_),
    .B1(_02274_),
    .B2(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__o22a_4 _16971_ (.A1(_06671_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02289_),
    .X(\CPU_src1_value_a2[19] ));
 sky130_fd_sc_hd__inv_2 _16972_ (.A(\CPU_Xreg_value_a4[8][20] ),
    .Y(_02290_));
 sky130_fd_sc_hd__a2bb2o_4 _16973_ (.A1_N(_02290_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][20] ),
    .B2(_02261_),
    .X(_02291_));
 sky130_fd_sc_hd__inv_2 _16974_ (.A(\CPU_Xreg_value_a4[5][20] ),
    .Y(_02292_));
 sky130_fd_sc_hd__inv_2 _16975_ (.A(\CPU_Xreg_value_a4[12][20] ),
    .Y(_02293_));
 sky130_fd_sc_hd__o22a_4 _16976_ (.A1(_02292_),
    .A2(_02221_),
    .B1(_02293_),
    .B2(_02223_),
    .X(_02294_));
 sky130_fd_sc_hd__inv_2 _16977_ (.A(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__inv_2 _16978_ (.A(\CPU_Xreg_value_a4[2][20] ),
    .Y(_02296_));
 sky130_fd_sc_hd__o21ai_4 _16979_ (.A1(_02296_),
    .A2(_02268_),
    .B1(_02194_),
    .Y(_02297_));
 sky130_fd_sc_hd__inv_2 _16980_ (.A(\CPU_Xreg_value_a4[14][20] ),
    .Y(_02298_));
 sky130_fd_sc_hd__inv_2 _16981_ (.A(\CPU_Xreg_value_a4[3][20] ),
    .Y(_02299_));
 sky130_fd_sc_hd__o22a_4 _16982_ (.A1(_02298_),
    .A2(_02229_),
    .B1(_02299_),
    .B2(_02231_),
    .X(_02300_));
 sky130_fd_sc_hd__inv_2 _16983_ (.A(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__or4_4 _16984_ (.A(_02291_),
    .B(_02295_),
    .C(_02297_),
    .D(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__inv_2 _16985_ (.A(\CPU_Xreg_value_a4[1][20] ),
    .Y(_02303_));
 sky130_fd_sc_hd__inv_2 _16986_ (.A(\CPU_Xreg_value_a4[4][20] ),
    .Y(_02304_));
 sky130_fd_sc_hd__o22a_4 _16987_ (.A1(_02303_),
    .A2(_02236_),
    .B1(_02304_),
    .B2(_02238_),
    .X(_02305_));
 sky130_fd_sc_hd__inv_2 _16988_ (.A(\CPU_Xreg_value_a4[6][20] ),
    .Y(_02306_));
 sky130_fd_sc_hd__inv_2 _16989_ (.A(\CPU_Xreg_value_a4[11][20] ),
    .Y(_02307_));
 sky130_fd_sc_hd__o22a_4 _16990_ (.A1(_02306_),
    .A2(_02241_),
    .B1(_02307_),
    .B2(_02243_),
    .X(_02308_));
 sky130_fd_sc_hd__inv_2 _16991_ (.A(\CPU_Xreg_value_a4[15][20] ),
    .Y(_02309_));
 sky130_fd_sc_hd__inv_2 _16992_ (.A(\CPU_Xreg_value_a4[10][20] ),
    .Y(_02310_));
 sky130_fd_sc_hd__o22a_4 _16993_ (.A1(_02309_),
    .A2(_02246_),
    .B1(_02310_),
    .B2(_02248_),
    .X(_02311_));
 sky130_fd_sc_hd__inv_2 _16994_ (.A(\CPU_Xreg_value_a4[9][20] ),
    .Y(_02312_));
 sky130_fd_sc_hd__inv_2 _16995_ (.A(\CPU_Xreg_value_a4[7][20] ),
    .Y(_02313_));
 sky130_fd_sc_hd__o22a_4 _16996_ (.A1(_02312_),
    .A2(_02251_),
    .B1(_02313_),
    .B2(_02253_),
    .X(_02314_));
 sky130_fd_sc_hd__and4_4 _16997_ (.A(_02305_),
    .B(_02308_),
    .C(_02311_),
    .D(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__inv_2 _16998_ (.A(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__o22a_4 _16999_ (.A1(\CPU_Xreg_value_a4[0][20] ),
    .A2(_02258_),
    .B1(_02302_),
    .B2(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__o22a_4 _17000_ (.A1(_06649_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02317_),
    .X(\CPU_src1_value_a2[20] ));
 sky130_fd_sc_hd__inv_2 _17001_ (.A(\CPU_Xreg_value_a4[8][21] ),
    .Y(_02318_));
 sky130_fd_sc_hd__a2bb2o_4 _17002_ (.A1_N(_02318_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][21] ),
    .B2(_02261_),
    .X(_02319_));
 sky130_fd_sc_hd__inv_2 _17003_ (.A(\CPU_Xreg_value_a4[5][21] ),
    .Y(_02320_));
 sky130_fd_sc_hd__inv_2 _17004_ (.A(\CPU_Xreg_value_a4[12][21] ),
    .Y(_02321_));
 sky130_fd_sc_hd__o22a_4 _17005_ (.A1(_02320_),
    .A2(_02221_),
    .B1(_02321_),
    .B2(_02223_),
    .X(_02322_));
 sky130_fd_sc_hd__inv_2 _17006_ (.A(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__inv_2 _17007_ (.A(\CPU_Xreg_value_a4[2][21] ),
    .Y(_02324_));
 sky130_fd_sc_hd__o21ai_4 _17008_ (.A1(_02324_),
    .A2(_02268_),
    .B1(_02194_),
    .Y(_02325_));
 sky130_fd_sc_hd__inv_2 _17009_ (.A(\CPU_Xreg_value_a4[14][21] ),
    .Y(_02326_));
 sky130_fd_sc_hd__inv_2 _17010_ (.A(\CPU_Xreg_value_a4[3][21] ),
    .Y(_02327_));
 sky130_fd_sc_hd__o22a_4 _17011_ (.A1(_02326_),
    .A2(_02229_),
    .B1(_02327_),
    .B2(_02231_),
    .X(_02328_));
 sky130_fd_sc_hd__inv_2 _17012_ (.A(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__or4_4 _17013_ (.A(_02319_),
    .B(_02323_),
    .C(_02325_),
    .D(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__inv_2 _17014_ (.A(\CPU_Xreg_value_a4[1][21] ),
    .Y(_02331_));
 sky130_fd_sc_hd__inv_2 _17015_ (.A(\CPU_Xreg_value_a4[4][21] ),
    .Y(_02332_));
 sky130_fd_sc_hd__o22a_4 _17016_ (.A1(_02331_),
    .A2(_02236_),
    .B1(_02332_),
    .B2(_02238_),
    .X(_02333_));
 sky130_fd_sc_hd__inv_2 _17017_ (.A(\CPU_Xreg_value_a4[6][21] ),
    .Y(_02334_));
 sky130_fd_sc_hd__inv_2 _17018_ (.A(\CPU_Xreg_value_a4[11][21] ),
    .Y(_02335_));
 sky130_fd_sc_hd__o22a_4 _17019_ (.A1(_02334_),
    .A2(_02241_),
    .B1(_02335_),
    .B2(_02243_),
    .X(_02336_));
 sky130_fd_sc_hd__inv_2 _17020_ (.A(\CPU_Xreg_value_a4[15][21] ),
    .Y(_02337_));
 sky130_fd_sc_hd__inv_2 _17021_ (.A(\CPU_Xreg_value_a4[10][21] ),
    .Y(_02338_));
 sky130_fd_sc_hd__o22a_4 _17022_ (.A1(_02337_),
    .A2(_02246_),
    .B1(_02338_),
    .B2(_02248_),
    .X(_02339_));
 sky130_fd_sc_hd__inv_2 _17023_ (.A(\CPU_Xreg_value_a4[9][21] ),
    .Y(_02340_));
 sky130_fd_sc_hd__inv_2 _17024_ (.A(\CPU_Xreg_value_a4[7][21] ),
    .Y(_02341_));
 sky130_fd_sc_hd__o22a_4 _17025_ (.A1(_02340_),
    .A2(_02251_),
    .B1(_02341_),
    .B2(_02253_),
    .X(_02342_));
 sky130_fd_sc_hd__and4_4 _17026_ (.A(_02333_),
    .B(_02336_),
    .C(_02339_),
    .D(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__inv_2 _17027_ (.A(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__o22a_4 _17028_ (.A1(\CPU_Xreg_value_a4[0][21] ),
    .A2(_02258_),
    .B1(_02330_),
    .B2(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__o22a_4 _17029_ (.A1(_06640_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02345_),
    .X(\CPU_src1_value_a2[21] ));
 sky130_fd_sc_hd__inv_2 _17030_ (.A(\CPU_Xreg_value_a4[8][22] ),
    .Y(_02346_));
 sky130_fd_sc_hd__a2bb2o_4 _17031_ (.A1_N(_02346_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][22] ),
    .B2(_02261_),
    .X(_02347_));
 sky130_fd_sc_hd__inv_2 _17032_ (.A(\CPU_Xreg_value_a4[5][22] ),
    .Y(_02348_));
 sky130_fd_sc_hd__inv_2 _17033_ (.A(\CPU_Xreg_value_a4[12][22] ),
    .Y(_02349_));
 sky130_fd_sc_hd__o22a_4 _17034_ (.A1(_02348_),
    .A2(_02221_),
    .B1(_02349_),
    .B2(_02223_),
    .X(_02350_));
 sky130_fd_sc_hd__inv_2 _17035_ (.A(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__inv_2 _17036_ (.A(\CPU_Xreg_value_a4[2][22] ),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_4 _17037_ (.A1(_02352_),
    .A2(_02268_),
    .B1(_02194_),
    .Y(_02353_));
 sky130_fd_sc_hd__inv_2 _17038_ (.A(\CPU_Xreg_value_a4[14][22] ),
    .Y(_02354_));
 sky130_fd_sc_hd__inv_2 _17039_ (.A(\CPU_Xreg_value_a4[3][22] ),
    .Y(_02355_));
 sky130_fd_sc_hd__o22a_4 _17040_ (.A1(_02354_),
    .A2(_02229_),
    .B1(_02355_),
    .B2(_02231_),
    .X(_02356_));
 sky130_fd_sc_hd__inv_2 _17041_ (.A(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__or4_4 _17042_ (.A(_02347_),
    .B(_02351_),
    .C(_02353_),
    .D(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__inv_2 _17043_ (.A(\CPU_Xreg_value_a4[1][22] ),
    .Y(_02359_));
 sky130_fd_sc_hd__inv_2 _17044_ (.A(\CPU_Xreg_value_a4[4][22] ),
    .Y(_02360_));
 sky130_fd_sc_hd__o22a_4 _17045_ (.A1(_02359_),
    .A2(_02236_),
    .B1(_02360_),
    .B2(_02238_),
    .X(_02361_));
 sky130_fd_sc_hd__inv_2 _17046_ (.A(\CPU_Xreg_value_a4[6][22] ),
    .Y(_02362_));
 sky130_fd_sc_hd__inv_2 _17047_ (.A(\CPU_Xreg_value_a4[11][22] ),
    .Y(_02363_));
 sky130_fd_sc_hd__o22a_4 _17048_ (.A1(_02362_),
    .A2(_02241_),
    .B1(_02363_),
    .B2(_02243_),
    .X(_02364_));
 sky130_fd_sc_hd__inv_2 _17049_ (.A(\CPU_Xreg_value_a4[15][22] ),
    .Y(_02365_));
 sky130_fd_sc_hd__inv_2 _17050_ (.A(\CPU_Xreg_value_a4[10][22] ),
    .Y(_02366_));
 sky130_fd_sc_hd__o22a_4 _17051_ (.A1(_02365_),
    .A2(_02246_),
    .B1(_02366_),
    .B2(_02248_),
    .X(_02367_));
 sky130_fd_sc_hd__inv_2 _17052_ (.A(\CPU_Xreg_value_a4[9][22] ),
    .Y(_02368_));
 sky130_fd_sc_hd__inv_2 _17053_ (.A(\CPU_Xreg_value_a4[7][22] ),
    .Y(_02369_));
 sky130_fd_sc_hd__o22a_4 _17054_ (.A1(_02368_),
    .A2(_02251_),
    .B1(_02369_),
    .B2(_02253_),
    .X(_02370_));
 sky130_fd_sc_hd__and4_4 _17055_ (.A(_02361_),
    .B(_02364_),
    .C(_02367_),
    .D(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__inv_2 _17056_ (.A(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o22a_4 _17057_ (.A1(\CPU_Xreg_value_a4[0][22] ),
    .A2(_02258_),
    .B1(_02358_),
    .B2(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__o22a_4 _17058_ (.A1(_06625_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02373_),
    .X(\CPU_src1_value_a2[22] ));
 sky130_fd_sc_hd__inv_2 _17059_ (.A(\CPU_Xreg_value_a4[8][23] ),
    .Y(_02374_));
 sky130_fd_sc_hd__a2bb2o_4 _17060_ (.A1_N(_02374_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][23] ),
    .B2(_02261_),
    .X(_02375_));
 sky130_fd_sc_hd__inv_2 _17061_ (.A(\CPU_Xreg_value_a4[5][23] ),
    .Y(_02376_));
 sky130_fd_sc_hd__inv_2 _17062_ (.A(\CPU_Xreg_value_a4[12][23] ),
    .Y(_02377_));
 sky130_fd_sc_hd__o22a_4 _17063_ (.A1(_02376_),
    .A2(_02221_),
    .B1(_02377_),
    .B2(_02223_),
    .X(_02378_));
 sky130_fd_sc_hd__inv_2 _17064_ (.A(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__inv_2 _17065_ (.A(\CPU_Xreg_value_a4[2][23] ),
    .Y(_02380_));
 sky130_fd_sc_hd__buf_2 _17066_ (.A(_01650_),
    .X(_02381_));
 sky130_fd_sc_hd__o21ai_4 _17067_ (.A1(_02380_),
    .A2(_02268_),
    .B1(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__inv_2 _17068_ (.A(\CPU_Xreg_value_a4[14][23] ),
    .Y(_02383_));
 sky130_fd_sc_hd__inv_2 _17069_ (.A(\CPU_Xreg_value_a4[3][23] ),
    .Y(_02384_));
 sky130_fd_sc_hd__o22a_4 _17070_ (.A1(_02383_),
    .A2(_02229_),
    .B1(_02384_),
    .B2(_02231_),
    .X(_02385_));
 sky130_fd_sc_hd__inv_2 _17071_ (.A(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__or4_4 _17072_ (.A(_02375_),
    .B(_02379_),
    .C(_02382_),
    .D(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__inv_2 _17073_ (.A(\CPU_Xreg_value_a4[1][23] ),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _17074_ (.A(\CPU_Xreg_value_a4[4][23] ),
    .Y(_02389_));
 sky130_fd_sc_hd__o22a_4 _17075_ (.A1(_02388_),
    .A2(_02236_),
    .B1(_02389_),
    .B2(_02238_),
    .X(_02390_));
 sky130_fd_sc_hd__inv_2 _17076_ (.A(\CPU_Xreg_value_a4[6][23] ),
    .Y(_02391_));
 sky130_fd_sc_hd__inv_2 _17077_ (.A(\CPU_Xreg_value_a4[11][23] ),
    .Y(_02392_));
 sky130_fd_sc_hd__o22a_4 _17078_ (.A1(_02391_),
    .A2(_02241_),
    .B1(_02392_),
    .B2(_02243_),
    .X(_02393_));
 sky130_fd_sc_hd__inv_2 _17079_ (.A(\CPU_Xreg_value_a4[15][23] ),
    .Y(_02394_));
 sky130_fd_sc_hd__inv_2 _17080_ (.A(\CPU_Xreg_value_a4[10][23] ),
    .Y(_02395_));
 sky130_fd_sc_hd__o22a_4 _17081_ (.A1(_02394_),
    .A2(_02246_),
    .B1(_02395_),
    .B2(_02248_),
    .X(_02396_));
 sky130_fd_sc_hd__inv_2 _17082_ (.A(\CPU_Xreg_value_a4[9][23] ),
    .Y(_02397_));
 sky130_fd_sc_hd__inv_2 _17083_ (.A(\CPU_Xreg_value_a4[7][23] ),
    .Y(_02398_));
 sky130_fd_sc_hd__o22a_4 _17084_ (.A1(_02397_),
    .A2(_02251_),
    .B1(_02398_),
    .B2(_02253_),
    .X(_02399_));
 sky130_fd_sc_hd__and4_4 _17085_ (.A(_02390_),
    .B(_02393_),
    .C(_02396_),
    .D(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__inv_2 _17086_ (.A(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__o22a_4 _17087_ (.A1(\CPU_Xreg_value_a4[0][23] ),
    .A2(_02258_),
    .B1(_02387_),
    .B2(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__o22a_4 _17088_ (.A1(_06617_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_02402_),
    .X(\CPU_src1_value_a2[23] ));
 sky130_fd_sc_hd__buf_2 _17089_ (.A(_01643_),
    .X(_02403_));
 sky130_fd_sc_hd__buf_2 _17090_ (.A(_01646_),
    .X(_02404_));
 sky130_fd_sc_hd__inv_2 _17091_ (.A(\CPU_Xreg_value_a4[8][24] ),
    .Y(_02405_));
 sky130_fd_sc_hd__a2bb2o_4 _17092_ (.A1_N(_02405_),
    .A2_N(_02260_),
    .B1(\CPU_Xreg_value_a4[13][24] ),
    .B2(_02261_),
    .X(_02406_));
 sky130_fd_sc_hd__inv_2 _17093_ (.A(\CPU_Xreg_value_a4[5][24] ),
    .Y(_02407_));
 sky130_fd_sc_hd__buf_2 _17094_ (.A(_01663_),
    .X(_02408_));
 sky130_fd_sc_hd__inv_2 _17095_ (.A(\CPU_Xreg_value_a4[12][24] ),
    .Y(_02409_));
 sky130_fd_sc_hd__buf_2 _17096_ (.A(_01667_),
    .X(_02410_));
 sky130_fd_sc_hd__o22a_4 _17097_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02409_),
    .B2(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__inv_2 _17098_ (.A(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _17099_ (.A(\CPU_Xreg_value_a4[2][24] ),
    .Y(_02413_));
 sky130_fd_sc_hd__o21ai_4 _17100_ (.A1(_02413_),
    .A2(_02268_),
    .B1(_02381_),
    .Y(_02414_));
 sky130_fd_sc_hd__inv_2 _17101_ (.A(\CPU_Xreg_value_a4[14][24] ),
    .Y(_02415_));
 sky130_fd_sc_hd__buf_2 _17102_ (.A(_01676_),
    .X(_02416_));
 sky130_fd_sc_hd__inv_2 _17103_ (.A(\CPU_Xreg_value_a4[3][24] ),
    .Y(_02417_));
 sky130_fd_sc_hd__buf_2 _17104_ (.A(_01679_),
    .X(_02418_));
 sky130_fd_sc_hd__o22a_4 _17105_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02417_),
    .B2(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__inv_2 _17106_ (.A(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__or4_4 _17107_ (.A(_02406_),
    .B(_02412_),
    .C(_02414_),
    .D(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__inv_2 _17108_ (.A(\CPU_Xreg_value_a4[1][24] ),
    .Y(_02422_));
 sky130_fd_sc_hd__buf_2 _17109_ (.A(_01684_),
    .X(_02423_));
 sky130_fd_sc_hd__inv_2 _17110_ (.A(\CPU_Xreg_value_a4[4][24] ),
    .Y(_02424_));
 sky130_fd_sc_hd__buf_2 _17111_ (.A(_01688_),
    .X(_02425_));
 sky130_fd_sc_hd__o22a_4 _17112_ (.A1(_02422_),
    .A2(_02423_),
    .B1(_02424_),
    .B2(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__inv_2 _17113_ (.A(\CPU_Xreg_value_a4[6][24] ),
    .Y(_02427_));
 sky130_fd_sc_hd__buf_2 _17114_ (.A(_01693_),
    .X(_02428_));
 sky130_fd_sc_hd__inv_2 _17115_ (.A(\CPU_Xreg_value_a4[11][24] ),
    .Y(_02429_));
 sky130_fd_sc_hd__buf_2 _17116_ (.A(_01696_),
    .X(_02430_));
 sky130_fd_sc_hd__o22a_4 _17117_ (.A1(_02427_),
    .A2(_02428_),
    .B1(_02429_),
    .B2(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__inv_2 _17118_ (.A(\CPU_Xreg_value_a4[15][24] ),
    .Y(_02432_));
 sky130_fd_sc_hd__buf_2 _17119_ (.A(_01700_),
    .X(_02433_));
 sky130_fd_sc_hd__inv_2 _17120_ (.A(\CPU_Xreg_value_a4[10][24] ),
    .Y(_02434_));
 sky130_fd_sc_hd__buf_2 _17121_ (.A(_01704_),
    .X(_02435_));
 sky130_fd_sc_hd__o22a_4 _17122_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02434_),
    .B2(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__inv_2 _17123_ (.A(\CPU_Xreg_value_a4[9][24] ),
    .Y(_02437_));
 sky130_fd_sc_hd__buf_2 _17124_ (.A(_01708_),
    .X(_02438_));
 sky130_fd_sc_hd__inv_2 _17125_ (.A(\CPU_Xreg_value_a4[7][24] ),
    .Y(_02439_));
 sky130_fd_sc_hd__buf_2 _17126_ (.A(_01711_),
    .X(_02440_));
 sky130_fd_sc_hd__o22a_4 _17127_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_02439_),
    .B2(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__and4_4 _17128_ (.A(_02426_),
    .B(_02431_),
    .C(_02436_),
    .D(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__inv_2 _17129_ (.A(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__o22a_4 _17130_ (.A1(\CPU_Xreg_value_a4[0][24] ),
    .A2(_02258_),
    .B1(_02421_),
    .B2(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__o22a_4 _17131_ (.A1(_06597_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02444_),
    .X(\CPU_src1_value_a2[24] ));
 sky130_fd_sc_hd__buf_2 _17132_ (.A(_01652_),
    .X(_02445_));
 sky130_fd_sc_hd__inv_2 _17133_ (.A(\CPU_Xreg_value_a4[8][25] ),
    .Y(_02446_));
 sky130_fd_sc_hd__buf_2 _17134_ (.A(_01656_),
    .X(_02447_));
 sky130_fd_sc_hd__buf_2 _17135_ (.A(_01721_),
    .X(_02448_));
 sky130_fd_sc_hd__a2bb2o_4 _17136_ (.A1_N(_02446_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][25] ),
    .B2(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__inv_2 _17137_ (.A(\CPU_Xreg_value_a4[5][25] ),
    .Y(_02450_));
 sky130_fd_sc_hd__inv_2 _17138_ (.A(\CPU_Xreg_value_a4[12][25] ),
    .Y(_02451_));
 sky130_fd_sc_hd__o22a_4 _17139_ (.A1(_02450_),
    .A2(_02408_),
    .B1(_02451_),
    .B2(_02410_),
    .X(_02452_));
 sky130_fd_sc_hd__inv_2 _17140_ (.A(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__inv_2 _17141_ (.A(\CPU_Xreg_value_a4[2][25] ),
    .Y(_02454_));
 sky130_fd_sc_hd__buf_2 _17142_ (.A(_01672_),
    .X(_02455_));
 sky130_fd_sc_hd__o21ai_4 _17143_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02381_),
    .Y(_02456_));
 sky130_fd_sc_hd__inv_2 _17144_ (.A(\CPU_Xreg_value_a4[14][25] ),
    .Y(_02457_));
 sky130_fd_sc_hd__inv_2 _17145_ (.A(\CPU_Xreg_value_a4[3][25] ),
    .Y(_02458_));
 sky130_fd_sc_hd__o22a_4 _17146_ (.A1(_02457_),
    .A2(_02416_),
    .B1(_02458_),
    .B2(_02418_),
    .X(_02459_));
 sky130_fd_sc_hd__inv_2 _17147_ (.A(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__or4_4 _17148_ (.A(_02449_),
    .B(_02453_),
    .C(_02456_),
    .D(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__inv_2 _17149_ (.A(\CPU_Xreg_value_a4[1][25] ),
    .Y(_02462_));
 sky130_fd_sc_hd__inv_2 _17150_ (.A(\CPU_Xreg_value_a4[4][25] ),
    .Y(_02463_));
 sky130_fd_sc_hd__o22a_4 _17151_ (.A1(_02462_),
    .A2(_02423_),
    .B1(_02463_),
    .B2(_02425_),
    .X(_02464_));
 sky130_fd_sc_hd__inv_2 _17152_ (.A(\CPU_Xreg_value_a4[6][25] ),
    .Y(_02465_));
 sky130_fd_sc_hd__inv_2 _17153_ (.A(\CPU_Xreg_value_a4[11][25] ),
    .Y(_02466_));
 sky130_fd_sc_hd__o22a_4 _17154_ (.A1(_02465_),
    .A2(_02428_),
    .B1(_02466_),
    .B2(_02430_),
    .X(_02467_));
 sky130_fd_sc_hd__inv_2 _17155_ (.A(\CPU_Xreg_value_a4[15][25] ),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _17156_ (.A(\CPU_Xreg_value_a4[10][25] ),
    .Y(_02469_));
 sky130_fd_sc_hd__o22a_4 _17157_ (.A1(_02468_),
    .A2(_02433_),
    .B1(_02469_),
    .B2(_02435_),
    .X(_02470_));
 sky130_fd_sc_hd__inv_2 _17158_ (.A(\CPU_Xreg_value_a4[9][25] ),
    .Y(_02471_));
 sky130_fd_sc_hd__inv_2 _17159_ (.A(\CPU_Xreg_value_a4[7][25] ),
    .Y(_02472_));
 sky130_fd_sc_hd__o22a_4 _17160_ (.A1(_02471_),
    .A2(_02438_),
    .B1(_02472_),
    .B2(_02440_),
    .X(_02473_));
 sky130_fd_sc_hd__and4_4 _17161_ (.A(_02464_),
    .B(_02467_),
    .C(_02470_),
    .D(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__inv_2 _17162_ (.A(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__o22a_4 _17163_ (.A1(\CPU_Xreg_value_a4[0][25] ),
    .A2(_02445_),
    .B1(_02461_),
    .B2(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__o22a_4 _17164_ (.A1(_06587_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02476_),
    .X(\CPU_src1_value_a2[25] ));
 sky130_fd_sc_hd__inv_2 _17165_ (.A(\CPU_Xreg_value_a4[8][26] ),
    .Y(_02477_));
 sky130_fd_sc_hd__a2bb2o_4 _17166_ (.A1_N(_02477_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][26] ),
    .B2(_02448_),
    .X(_02478_));
 sky130_fd_sc_hd__inv_2 _17167_ (.A(\CPU_Xreg_value_a4[5][26] ),
    .Y(_02479_));
 sky130_fd_sc_hd__inv_2 _17168_ (.A(\CPU_Xreg_value_a4[12][26] ),
    .Y(_02480_));
 sky130_fd_sc_hd__o22a_4 _17169_ (.A1(_02479_),
    .A2(_02408_),
    .B1(_02480_),
    .B2(_02410_),
    .X(_02481_));
 sky130_fd_sc_hd__inv_2 _17170_ (.A(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__inv_2 _17171_ (.A(\CPU_Xreg_value_a4[2][26] ),
    .Y(_02483_));
 sky130_fd_sc_hd__o21ai_4 _17172_ (.A1(_02483_),
    .A2(_02455_),
    .B1(_02381_),
    .Y(_02484_));
 sky130_fd_sc_hd__inv_2 _17173_ (.A(\CPU_Xreg_value_a4[14][26] ),
    .Y(_02485_));
 sky130_fd_sc_hd__inv_2 _17174_ (.A(\CPU_Xreg_value_a4[3][26] ),
    .Y(_02486_));
 sky130_fd_sc_hd__o22a_4 _17175_ (.A1(_02485_),
    .A2(_02416_),
    .B1(_02486_),
    .B2(_02418_),
    .X(_02487_));
 sky130_fd_sc_hd__inv_2 _17176_ (.A(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__or4_4 _17177_ (.A(_02478_),
    .B(_02482_),
    .C(_02484_),
    .D(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__inv_2 _17178_ (.A(\CPU_Xreg_value_a4[1][26] ),
    .Y(_02490_));
 sky130_fd_sc_hd__inv_2 _17179_ (.A(\CPU_Xreg_value_a4[4][26] ),
    .Y(_02491_));
 sky130_fd_sc_hd__o22a_4 _17180_ (.A1(_02490_),
    .A2(_02423_),
    .B1(_02491_),
    .B2(_02425_),
    .X(_02492_));
 sky130_fd_sc_hd__inv_2 _17181_ (.A(\CPU_Xreg_value_a4[6][26] ),
    .Y(_02493_));
 sky130_fd_sc_hd__inv_2 _17182_ (.A(\CPU_Xreg_value_a4[11][26] ),
    .Y(_02494_));
 sky130_fd_sc_hd__o22a_4 _17183_ (.A1(_02493_),
    .A2(_02428_),
    .B1(_02494_),
    .B2(_02430_),
    .X(_02495_));
 sky130_fd_sc_hd__inv_2 _17184_ (.A(\CPU_Xreg_value_a4[15][26] ),
    .Y(_02496_));
 sky130_fd_sc_hd__inv_2 _17185_ (.A(\CPU_Xreg_value_a4[10][26] ),
    .Y(_02497_));
 sky130_fd_sc_hd__o22a_4 _17186_ (.A1(_02496_),
    .A2(_02433_),
    .B1(_02497_),
    .B2(_02435_),
    .X(_02498_));
 sky130_fd_sc_hd__inv_2 _17187_ (.A(\CPU_Xreg_value_a4[9][26] ),
    .Y(_02499_));
 sky130_fd_sc_hd__inv_2 _17188_ (.A(\CPU_Xreg_value_a4[7][26] ),
    .Y(_02500_));
 sky130_fd_sc_hd__o22a_4 _17189_ (.A1(_02499_),
    .A2(_02438_),
    .B1(_02500_),
    .B2(_02440_),
    .X(_02501_));
 sky130_fd_sc_hd__and4_4 _17190_ (.A(_02492_),
    .B(_02495_),
    .C(_02498_),
    .D(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__inv_2 _17191_ (.A(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__o22a_4 _17192_ (.A1(\CPU_Xreg_value_a4[0][26] ),
    .A2(_02445_),
    .B1(_02489_),
    .B2(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__o22a_4 _17193_ (.A1(_06572_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02504_),
    .X(\CPU_src1_value_a2[26] ));
 sky130_fd_sc_hd__inv_2 _17194_ (.A(\CPU_Xreg_value_a4[8][27] ),
    .Y(_02505_));
 sky130_fd_sc_hd__a2bb2o_4 _17195_ (.A1_N(_02505_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][27] ),
    .B2(_02448_),
    .X(_02506_));
 sky130_fd_sc_hd__inv_2 _17196_ (.A(\CPU_Xreg_value_a4[5][27] ),
    .Y(_02507_));
 sky130_fd_sc_hd__inv_2 _17197_ (.A(\CPU_Xreg_value_a4[12][27] ),
    .Y(_02508_));
 sky130_fd_sc_hd__o22a_4 _17198_ (.A1(_02507_),
    .A2(_02408_),
    .B1(_02508_),
    .B2(_02410_),
    .X(_02509_));
 sky130_fd_sc_hd__inv_2 _17199_ (.A(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _17200_ (.A(\CPU_Xreg_value_a4[2][27] ),
    .Y(_02511_));
 sky130_fd_sc_hd__o21ai_4 _17201_ (.A1(_02511_),
    .A2(_02455_),
    .B1(_02381_),
    .Y(_02512_));
 sky130_fd_sc_hd__inv_2 _17202_ (.A(\CPU_Xreg_value_a4[14][27] ),
    .Y(_02513_));
 sky130_fd_sc_hd__inv_2 _17203_ (.A(\CPU_Xreg_value_a4[3][27] ),
    .Y(_02514_));
 sky130_fd_sc_hd__o22a_4 _17204_ (.A1(_02513_),
    .A2(_02416_),
    .B1(_02514_),
    .B2(_02418_),
    .X(_02515_));
 sky130_fd_sc_hd__inv_2 _17205_ (.A(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__or4_4 _17206_ (.A(_02506_),
    .B(_02510_),
    .C(_02512_),
    .D(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__inv_2 _17207_ (.A(\CPU_Xreg_value_a4[1][27] ),
    .Y(_02518_));
 sky130_fd_sc_hd__inv_2 _17208_ (.A(\CPU_Xreg_value_a4[4][27] ),
    .Y(_02519_));
 sky130_fd_sc_hd__o22a_4 _17209_ (.A1(_02518_),
    .A2(_02423_),
    .B1(_02519_),
    .B2(_02425_),
    .X(_02520_));
 sky130_fd_sc_hd__inv_2 _17210_ (.A(\CPU_Xreg_value_a4[6][27] ),
    .Y(_02521_));
 sky130_fd_sc_hd__inv_2 _17211_ (.A(\CPU_Xreg_value_a4[11][27] ),
    .Y(_02522_));
 sky130_fd_sc_hd__o22a_4 _17212_ (.A1(_02521_),
    .A2(_02428_),
    .B1(_02522_),
    .B2(_02430_),
    .X(_02523_));
 sky130_fd_sc_hd__inv_2 _17213_ (.A(\CPU_Xreg_value_a4[15][27] ),
    .Y(_02524_));
 sky130_fd_sc_hd__inv_2 _17214_ (.A(\CPU_Xreg_value_a4[10][27] ),
    .Y(_02525_));
 sky130_fd_sc_hd__o22a_4 _17215_ (.A1(_02524_),
    .A2(_02433_),
    .B1(_02525_),
    .B2(_02435_),
    .X(_02526_));
 sky130_fd_sc_hd__inv_2 _17216_ (.A(\CPU_Xreg_value_a4[9][27] ),
    .Y(_02527_));
 sky130_fd_sc_hd__inv_2 _17217_ (.A(\CPU_Xreg_value_a4[7][27] ),
    .Y(_02528_));
 sky130_fd_sc_hd__o22a_4 _17218_ (.A1(_02527_),
    .A2(_02438_),
    .B1(_02528_),
    .B2(_02440_),
    .X(_02529_));
 sky130_fd_sc_hd__and4_4 _17219_ (.A(_02520_),
    .B(_02523_),
    .C(_02526_),
    .D(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__inv_2 _17220_ (.A(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__o22a_4 _17221_ (.A1(\CPU_Xreg_value_a4[0][27] ),
    .A2(_02445_),
    .B1(_02517_),
    .B2(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__o22a_4 _17222_ (.A1(_06562_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02532_),
    .X(\CPU_src1_value_a2[27] ));
 sky130_fd_sc_hd__inv_2 _17223_ (.A(\CPU_Xreg_value_a4[8][28] ),
    .Y(_02533_));
 sky130_fd_sc_hd__a2bb2o_4 _17224_ (.A1_N(_02533_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][28] ),
    .B2(_02448_),
    .X(_02534_));
 sky130_fd_sc_hd__inv_2 _17225_ (.A(\CPU_Xreg_value_a4[5][28] ),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_2 _17226_ (.A(\CPU_Xreg_value_a4[12][28] ),
    .Y(_02536_));
 sky130_fd_sc_hd__o22a_4 _17227_ (.A1(_02535_),
    .A2(_02408_),
    .B1(_02536_),
    .B2(_02410_),
    .X(_02537_));
 sky130_fd_sc_hd__inv_2 _17228_ (.A(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__inv_2 _17229_ (.A(\CPU_Xreg_value_a4[2][28] ),
    .Y(_02539_));
 sky130_fd_sc_hd__o21ai_4 _17230_ (.A1(_02539_),
    .A2(_02455_),
    .B1(_02381_),
    .Y(_02540_));
 sky130_fd_sc_hd__inv_2 _17231_ (.A(\CPU_Xreg_value_a4[14][28] ),
    .Y(_02541_));
 sky130_fd_sc_hd__inv_2 _17232_ (.A(\CPU_Xreg_value_a4[3][28] ),
    .Y(_02542_));
 sky130_fd_sc_hd__o22a_4 _17233_ (.A1(_02541_),
    .A2(_02416_),
    .B1(_02542_),
    .B2(_02418_),
    .X(_02543_));
 sky130_fd_sc_hd__inv_2 _17234_ (.A(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__or4_4 _17235_ (.A(_02534_),
    .B(_02538_),
    .C(_02540_),
    .D(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__inv_2 _17236_ (.A(\CPU_Xreg_value_a4[1][28] ),
    .Y(_02546_));
 sky130_fd_sc_hd__inv_2 _17237_ (.A(\CPU_Xreg_value_a4[4][28] ),
    .Y(_02547_));
 sky130_fd_sc_hd__o22a_4 _17238_ (.A1(_02546_),
    .A2(_02423_),
    .B1(_02547_),
    .B2(_02425_),
    .X(_02548_));
 sky130_fd_sc_hd__inv_2 _17239_ (.A(\CPU_Xreg_value_a4[6][28] ),
    .Y(_02549_));
 sky130_fd_sc_hd__inv_2 _17240_ (.A(\CPU_Xreg_value_a4[11][28] ),
    .Y(_02550_));
 sky130_fd_sc_hd__o22a_4 _17241_ (.A1(_02549_),
    .A2(_02428_),
    .B1(_02550_),
    .B2(_02430_),
    .X(_02551_));
 sky130_fd_sc_hd__inv_2 _17242_ (.A(\CPU_Xreg_value_a4[15][28] ),
    .Y(_02552_));
 sky130_fd_sc_hd__inv_2 _17243_ (.A(\CPU_Xreg_value_a4[10][28] ),
    .Y(_02553_));
 sky130_fd_sc_hd__o22a_4 _17244_ (.A1(_02552_),
    .A2(_02433_),
    .B1(_02553_),
    .B2(_02435_),
    .X(_02554_));
 sky130_fd_sc_hd__inv_2 _17245_ (.A(\CPU_Xreg_value_a4[9][28] ),
    .Y(_02555_));
 sky130_fd_sc_hd__inv_2 _17246_ (.A(\CPU_Xreg_value_a4[7][28] ),
    .Y(_02556_));
 sky130_fd_sc_hd__o22a_4 _17247_ (.A1(_02555_),
    .A2(_02438_),
    .B1(_02556_),
    .B2(_02440_),
    .X(_02557_));
 sky130_fd_sc_hd__and4_4 _17248_ (.A(_02548_),
    .B(_02551_),
    .C(_02554_),
    .D(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__inv_2 _17249_ (.A(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__o22a_4 _17250_ (.A1(\CPU_Xreg_value_a4[0][28] ),
    .A2(_02445_),
    .B1(_02545_),
    .B2(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__o22a_4 _17251_ (.A1(_06537_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02560_),
    .X(\CPU_src1_value_a2[28] ));
 sky130_fd_sc_hd__inv_2 _17252_ (.A(\CPU_Xreg_value_a4[8][29] ),
    .Y(_02561_));
 sky130_fd_sc_hd__a2bb2o_4 _17253_ (.A1_N(_02561_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][29] ),
    .B2(_02448_),
    .X(_02562_));
 sky130_fd_sc_hd__inv_2 _17254_ (.A(\CPU_Xreg_value_a4[5][29] ),
    .Y(_02563_));
 sky130_fd_sc_hd__inv_2 _17255_ (.A(\CPU_Xreg_value_a4[12][29] ),
    .Y(_02564_));
 sky130_fd_sc_hd__o22a_4 _17256_ (.A1(_02563_),
    .A2(_02408_),
    .B1(_02564_),
    .B2(_02410_),
    .X(_02565_));
 sky130_fd_sc_hd__inv_2 _17257_ (.A(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__inv_2 _17258_ (.A(\CPU_Xreg_value_a4[2][29] ),
    .Y(_02567_));
 sky130_fd_sc_hd__o21ai_4 _17259_ (.A1(_02567_),
    .A2(_02455_),
    .B1(_01651_),
    .Y(_02568_));
 sky130_fd_sc_hd__inv_2 _17260_ (.A(\CPU_Xreg_value_a4[14][29] ),
    .Y(_02569_));
 sky130_fd_sc_hd__inv_2 _17261_ (.A(\CPU_Xreg_value_a4[3][29] ),
    .Y(_02570_));
 sky130_fd_sc_hd__o22a_4 _17262_ (.A1(_02569_),
    .A2(_02416_),
    .B1(_02570_),
    .B2(_02418_),
    .X(_02571_));
 sky130_fd_sc_hd__inv_2 _17263_ (.A(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__or4_4 _17264_ (.A(_02562_),
    .B(_02566_),
    .C(_02568_),
    .D(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__inv_2 _17265_ (.A(\CPU_Xreg_value_a4[1][29] ),
    .Y(_02574_));
 sky130_fd_sc_hd__inv_2 _17266_ (.A(\CPU_Xreg_value_a4[4][29] ),
    .Y(_02575_));
 sky130_fd_sc_hd__o22a_4 _17267_ (.A1(_02574_),
    .A2(_02423_),
    .B1(_02575_),
    .B2(_02425_),
    .X(_02576_));
 sky130_fd_sc_hd__inv_2 _17268_ (.A(\CPU_Xreg_value_a4[6][29] ),
    .Y(_02577_));
 sky130_fd_sc_hd__inv_2 _17269_ (.A(\CPU_Xreg_value_a4[11][29] ),
    .Y(_02578_));
 sky130_fd_sc_hd__o22a_4 _17270_ (.A1(_02577_),
    .A2(_02428_),
    .B1(_02578_),
    .B2(_02430_),
    .X(_02579_));
 sky130_fd_sc_hd__inv_2 _17271_ (.A(\CPU_Xreg_value_a4[15][29] ),
    .Y(_02580_));
 sky130_fd_sc_hd__inv_2 _17272_ (.A(\CPU_Xreg_value_a4[10][29] ),
    .Y(_02581_));
 sky130_fd_sc_hd__o22a_4 _17273_ (.A1(_02580_),
    .A2(_02433_),
    .B1(_02581_),
    .B2(_02435_),
    .X(_02582_));
 sky130_fd_sc_hd__inv_2 _17274_ (.A(\CPU_Xreg_value_a4[9][29] ),
    .Y(_02583_));
 sky130_fd_sc_hd__inv_2 _17275_ (.A(\CPU_Xreg_value_a4[7][29] ),
    .Y(_02584_));
 sky130_fd_sc_hd__o22a_4 _17276_ (.A1(_02583_),
    .A2(_02438_),
    .B1(_02584_),
    .B2(_02440_),
    .X(_02585_));
 sky130_fd_sc_hd__and4_4 _17277_ (.A(_02576_),
    .B(_02579_),
    .C(_02582_),
    .D(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__inv_2 _17278_ (.A(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__o22a_4 _17279_ (.A1(\CPU_Xreg_value_a4[0][29] ),
    .A2(_02445_),
    .B1(_02573_),
    .B2(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__o22a_4 _17280_ (.A1(_06529_),
    .A2(_02403_),
    .B1(_02404_),
    .B2(_02588_),
    .X(\CPU_src1_value_a2[29] ));
 sky130_fd_sc_hd__inv_2 _17281_ (.A(\CPU_Xreg_value_a4[8][30] ),
    .Y(_02589_));
 sky130_fd_sc_hd__a2bb2o_4 _17282_ (.A1_N(_02589_),
    .A2_N(_02447_),
    .B1(\CPU_Xreg_value_a4[13][30] ),
    .B2(_02448_),
    .X(_02590_));
 sky130_fd_sc_hd__inv_2 _17283_ (.A(\CPU_Xreg_value_a4[5][30] ),
    .Y(_02591_));
 sky130_fd_sc_hd__inv_2 _17284_ (.A(\CPU_Xreg_value_a4[12][30] ),
    .Y(_02592_));
 sky130_fd_sc_hd__o22a_4 _17285_ (.A1(_02591_),
    .A2(_01664_),
    .B1(_02592_),
    .B2(_01668_),
    .X(_02593_));
 sky130_fd_sc_hd__inv_2 _17286_ (.A(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__inv_2 _17287_ (.A(\CPU_Xreg_value_a4[2][30] ),
    .Y(_02595_));
 sky130_fd_sc_hd__o21ai_4 _17288_ (.A1(_02595_),
    .A2(_02455_),
    .B1(_01651_),
    .Y(_02596_));
 sky130_fd_sc_hd__inv_2 _17289_ (.A(\CPU_Xreg_value_a4[14][30] ),
    .Y(_02597_));
 sky130_fd_sc_hd__inv_2 _17290_ (.A(\CPU_Xreg_value_a4[3][30] ),
    .Y(_02598_));
 sky130_fd_sc_hd__o22a_4 _17291_ (.A1(_02597_),
    .A2(_01677_),
    .B1(_02598_),
    .B2(_01680_),
    .X(_02599_));
 sky130_fd_sc_hd__inv_2 _17292_ (.A(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__or4_4 _17293_ (.A(_02590_),
    .B(_02594_),
    .C(_02596_),
    .D(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__inv_2 _17294_ (.A(\CPU_Xreg_value_a4[1][30] ),
    .Y(_02602_));
 sky130_fd_sc_hd__inv_2 _17295_ (.A(\CPU_Xreg_value_a4[4][30] ),
    .Y(_02603_));
 sky130_fd_sc_hd__o22a_4 _17296_ (.A1(_02602_),
    .A2(_01685_),
    .B1(_02603_),
    .B2(_01689_),
    .X(_02604_));
 sky130_fd_sc_hd__inv_2 _17297_ (.A(\CPU_Xreg_value_a4[6][30] ),
    .Y(_02605_));
 sky130_fd_sc_hd__inv_2 _17298_ (.A(\CPU_Xreg_value_a4[11][30] ),
    .Y(_02606_));
 sky130_fd_sc_hd__o22a_4 _17299_ (.A1(_02605_),
    .A2(_01694_),
    .B1(_02606_),
    .B2(_01697_),
    .X(_02607_));
 sky130_fd_sc_hd__inv_2 _17300_ (.A(\CPU_Xreg_value_a4[15][30] ),
    .Y(_02608_));
 sky130_fd_sc_hd__inv_2 _17301_ (.A(\CPU_Xreg_value_a4[10][30] ),
    .Y(_02609_));
 sky130_fd_sc_hd__o22a_4 _17302_ (.A1(_02608_),
    .A2(_01701_),
    .B1(_02609_),
    .B2(_01705_),
    .X(_02610_));
 sky130_fd_sc_hd__inv_2 _17303_ (.A(\CPU_Xreg_value_a4[9][30] ),
    .Y(_02611_));
 sky130_fd_sc_hd__inv_2 _17304_ (.A(\CPU_Xreg_value_a4[7][30] ),
    .Y(_02612_));
 sky130_fd_sc_hd__o22a_4 _17305_ (.A1(_02611_),
    .A2(_01709_),
    .B1(_02612_),
    .B2(_01712_),
    .X(_02613_));
 sky130_fd_sc_hd__and4_4 _17306_ (.A(_02604_),
    .B(_02607_),
    .C(_02610_),
    .D(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__inv_2 _17307_ (.A(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__o22a_4 _17308_ (.A1(\CPU_Xreg_value_a4[0][30] ),
    .A2(_02445_),
    .B1(_02601_),
    .B2(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__o22a_4 _17309_ (.A1(_06513_),
    .A2(_01644_),
    .B1(_01647_),
    .B2(_02616_),
    .X(\CPU_src1_value_a2[30] ));
 sky130_fd_sc_hd__inv_2 _17310_ (.A(\CPU_Xreg_value_a4[8][31] ),
    .Y(_02617_));
 sky130_fd_sc_hd__a2bb2o_4 _17311_ (.A1_N(_02617_),
    .A2_N(_01657_),
    .B1(\CPU_Xreg_value_a4[13][31] ),
    .B2(_01721_),
    .X(_02618_));
 sky130_fd_sc_hd__inv_2 _17312_ (.A(\CPU_Xreg_value_a4[5][31] ),
    .Y(_02619_));
 sky130_fd_sc_hd__inv_2 _17313_ (.A(\CPU_Xreg_value_a4[12][31] ),
    .Y(_02620_));
 sky130_fd_sc_hd__o22a_4 _17314_ (.A1(_02619_),
    .A2(_01664_),
    .B1(_02620_),
    .B2(_01668_),
    .X(_02621_));
 sky130_fd_sc_hd__inv_2 _17315_ (.A(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__inv_2 _17316_ (.A(\CPU_Xreg_value_a4[2][31] ),
    .Y(_02623_));
 sky130_fd_sc_hd__o21ai_4 _17317_ (.A1(_02623_),
    .A2(_01673_),
    .B1(_01651_),
    .Y(_02624_));
 sky130_fd_sc_hd__inv_2 _17318_ (.A(\CPU_Xreg_value_a4[14][31] ),
    .Y(_02625_));
 sky130_fd_sc_hd__inv_2 _17319_ (.A(\CPU_Xreg_value_a4[3][31] ),
    .Y(_02626_));
 sky130_fd_sc_hd__o22a_4 _17320_ (.A1(_02625_),
    .A2(_01677_),
    .B1(_02626_),
    .B2(_01680_),
    .X(_02627_));
 sky130_fd_sc_hd__inv_2 _17321_ (.A(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__or4_4 _17322_ (.A(_02618_),
    .B(_02622_),
    .C(_02624_),
    .D(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__inv_2 _17323_ (.A(\CPU_Xreg_value_a4[1][31] ),
    .Y(_02630_));
 sky130_fd_sc_hd__inv_2 _17324_ (.A(\CPU_Xreg_value_a4[4][31] ),
    .Y(_02631_));
 sky130_fd_sc_hd__o22a_4 _17325_ (.A1(_02630_),
    .A2(_01685_),
    .B1(_02631_),
    .B2(_01689_),
    .X(_02632_));
 sky130_fd_sc_hd__inv_2 _17326_ (.A(\CPU_Xreg_value_a4[6][31] ),
    .Y(_02633_));
 sky130_fd_sc_hd__inv_2 _17327_ (.A(\CPU_Xreg_value_a4[11][31] ),
    .Y(_02634_));
 sky130_fd_sc_hd__o22a_4 _17328_ (.A1(_02633_),
    .A2(_01694_),
    .B1(_02634_),
    .B2(_01697_),
    .X(_02635_));
 sky130_fd_sc_hd__inv_2 _17329_ (.A(\CPU_Xreg_value_a4[15][31] ),
    .Y(_02636_));
 sky130_fd_sc_hd__inv_2 _17330_ (.A(\CPU_Xreg_value_a4[10][31] ),
    .Y(_02637_));
 sky130_fd_sc_hd__o22a_4 _17331_ (.A1(_02636_),
    .A2(_01701_),
    .B1(_02637_),
    .B2(_01705_),
    .X(_02638_));
 sky130_fd_sc_hd__inv_2 _17332_ (.A(\CPU_Xreg_value_a4[9][31] ),
    .Y(_02639_));
 sky130_fd_sc_hd__inv_2 _17333_ (.A(\CPU_Xreg_value_a4[7][31] ),
    .Y(_02640_));
 sky130_fd_sc_hd__o22a_4 _17334_ (.A1(_02639_),
    .A2(_01709_),
    .B1(_02640_),
    .B2(_01712_),
    .X(_02641_));
 sky130_fd_sc_hd__and4_4 _17335_ (.A(_02632_),
    .B(_02635_),
    .C(_02638_),
    .D(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__inv_2 _17336_ (.A(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__o22a_4 _17337_ (.A1(\CPU_Xreg_value_a4[0][31] ),
    .A2(_01653_),
    .B1(_02629_),
    .B2(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__o22a_4 _17338_ (.A1(_06501_),
    .A2(_01644_),
    .B1(_01647_),
    .B2(_02644_),
    .X(\CPU_src1_value_a2[31] ));
 sky130_fd_sc_hd__inv_2 _17339_ (.A(\CPU_rf_rd_index2_a2[0] ),
    .Y(_02645_));
 sky130_fd_sc_hd__buf_2 _17340_ (.A(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__a2bb2o_4 _17341_ (.A1_N(\CPU_rd_a3[0] ),
    .A2_N(_02646_),
    .B1(\CPU_rd_a3[0] ),
    .B2(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__inv_2 _17342_ (.A(\CPU_rd_a3[1] ),
    .Y(_02648_));
 sky130_fd_sc_hd__buf_2 _17343_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .X(_02649_));
 sky130_fd_sc_hd__buf_2 _17344_ (.A(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__inv_2 _17345_ (.A(\CPU_rf_rd_index2_a2[4] ),
    .Y(_02651_));
 sky130_fd_sc_hd__buf_2 _17346_ (.A(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__buf_2 _17347_ (.A(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__o22a_4 _17348_ (.A1(_02648_),
    .A2(_02650_),
    .B1(\CPU_rd_a3[4] ),
    .B2(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__inv_2 _17349_ (.A(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__and2_4 _17350_ (.A(\CPU_rd_a3[4] ),
    .B(_02653_),
    .X(_02656_));
 sky130_fd_sc_hd__buf_2 _17351_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .X(_02657_));
 sky130_fd_sc_hd__buf_2 _17352_ (.A(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__buf_2 _17353_ (.A(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__a2bb2o_4 _17354_ (.A1_N(_01630_),
    .A2_N(_02659_),
    .B1(_01630_),
    .B2(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__buf_2 _17355_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .X(_02661_));
 sky130_fd_sc_hd__buf_2 _17356_ (.A(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__inv_2 _17357_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .Y(_02663_));
 sky130_fd_sc_hd__buf_2 _17358_ (.A(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__buf_2 _17359_ (.A(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__o22a_4 _17360_ (.A1(\CPU_rd_a3[3] ),
    .A2(_02662_),
    .B1(_01633_),
    .B2(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__a2111o_4 _17361_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_02656_),
    .C1(_02660_),
    .D1(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__or4_4 _17362_ (.A(_02647_),
    .B(_02655_),
    .C(_02667_),
    .D(_01642_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_2 _17363_ (.A(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__buf_2 _17364_ (.A(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__inv_2 _17365_ (.A(_02668_),
    .Y(_02671_));
 sky130_fd_sc_hd__buf_2 _17366_ (.A(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__buf_2 _17367_ (.A(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__inv_2 _17368_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .Y(_02674_));
 sky130_fd_sc_hd__or2_4 _17369_ (.A(_02674_),
    .B(_02645_),
    .X(_02675_));
 sky130_fd_sc_hd__buf_2 _17370_ (.A(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__buf_2 _17371_ (.A(\CPU_rf_rd_index2_a2[4] ),
    .X(_02677_));
 sky130_fd_sc_hd__buf_2 _17372_ (.A(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_2 _17373_ (.A(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__or4_4 _17374_ (.A(_02662_),
    .B(_02659_),
    .C(_02676_),
    .D(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__buf_2 _17375_ (.A(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__buf_2 _17376_ (.A(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__or2_4 _17377_ (.A(_02674_),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .X(_02683_));
 sky130_fd_sc_hd__buf_2 _17378_ (.A(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__or4_4 _17379_ (.A(_02665_),
    .B(_02659_),
    .C(_02684_),
    .D(_02679_),
    .X(_02685_));
 sky130_fd_sc_hd__buf_2 _17380_ (.A(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__buf_2 _17381_ (.A(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__o22a_4 _17382_ (.A1(_07189_),
    .A2(_02682_),
    .B1(_01703_),
    .B2(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__or2_4 _17383_ (.A(_02649_),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .X(_02689_));
 sky130_fd_sc_hd__buf_2 _17384_ (.A(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__or4_4 _17385_ (.A(_02661_),
    .B(_02658_),
    .C(_02690_),
    .D(_02652_),
    .X(_02691_));
 sky130_fd_sc_hd__inv_2 _17386_ (.A(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__buf_2 _17387_ (.A(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__buf_2 _17388_ (.A(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__inv_2 _17389_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .Y(_02695_));
 sky130_fd_sc_hd__buf_2 _17390_ (.A(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__or4_4 _17391_ (.A(_02664_),
    .B(_02696_),
    .C(_02684_),
    .D(_02653_),
    .X(_02697_));
 sky130_fd_sc_hd__inv_2 _17392_ (.A(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__buf_2 _17393_ (.A(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__buf_2 _17394_ (.A(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__a22oi_4 _17395_ (.A1(\CPU_Xreg_value_a4[16][0] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][0] ),
    .B2(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__buf_2 _17396_ (.A(_02696_),
    .X(_02702_));
 sky130_fd_sc_hd__or4_4 _17397_ (.A(_02662_),
    .B(_02702_),
    .C(_02684_),
    .D(_02678_),
    .X(_02703_));
 sky130_fd_sc_hd__buf_2 _17398_ (.A(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__buf_2 _17399_ (.A(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__or2_4 _17400_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .B(_02695_),
    .X(_02706_));
 sky130_fd_sc_hd__or4_4 _17401_ (.A(_02650_),
    .B(_02646_),
    .C(_02706_),
    .D(_02679_),
    .X(_02707_));
 sky130_fd_sc_hd__buf_2 _17402_ (.A(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__buf_2 _17403_ (.A(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__o22a_4 _17404_ (.A1(_01692_),
    .A2(_02705_),
    .B1(_07363_),
    .B2(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__or4_4 _17405_ (.A(_02662_),
    .B(_02702_),
    .C(_02690_),
    .D(_02678_),
    .X(_02711_));
 sky130_fd_sc_hd__buf_2 _17406_ (.A(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__buf_2 _17407_ (.A(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__or4_4 _17408_ (.A(_02665_),
    .B(_02659_),
    .C(_02676_),
    .D(_02679_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_2 _17409_ (.A(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__buf_2 _17410_ (.A(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__o22a_4 _17411_ (.A1(_01687_),
    .A2(_02713_),
    .B1(_07902_),
    .B2(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__and4_4 _17412_ (.A(_02688_),
    .B(_02701_),
    .C(_02710_),
    .D(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__inv_2 _17413_ (.A(\CPU_Xreg_value_a4[26][0] ),
    .Y(_02719_));
 sky130_fd_sc_hd__or4_4 _17414_ (.A(_02665_),
    .B(_02659_),
    .C(_02684_),
    .D(_02653_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_2 _17415_ (.A(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__buf_2 _17416_ (.A(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__or4_4 _17417_ (.A(_02665_),
    .B(_02702_),
    .C(_02690_),
    .D(_02679_),
    .X(_02723_));
 sky130_fd_sc_hd__buf_2 _17418_ (.A(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__buf_2 _17419_ (.A(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__o22a_4 _17420_ (.A1(_02719_),
    .A2(_02722_),
    .B1(_01666_),
    .B2(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__or4_4 _17421_ (.A(_02664_),
    .B(_02702_),
    .C(_02676_),
    .D(_02678_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_2 _17422_ (.A(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__buf_2 _17423_ (.A(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__or4_4 _17424_ (.A(_02665_),
    .B(_02702_),
    .C(_02684_),
    .D(_02679_),
    .X(_02730_));
 sky130_fd_sc_hd__buf_2 _17425_ (.A(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__buf_2 _17426_ (.A(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__o22a_4 _17427_ (.A1(_08271_),
    .A2(_02729_),
    .B1(_01675_),
    .B2(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__or4_4 _17428_ (.A(_02661_),
    .B(_02696_),
    .C(_02675_),
    .D(_02652_),
    .X(_02734_));
 sky130_fd_sc_hd__inv_2 _17429_ (.A(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__buf_2 _17430_ (.A(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__buf_2 _17431_ (.A(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__or4_4 _17432_ (.A(_02664_),
    .B(_02696_),
    .C(_02676_),
    .D(_02653_),
    .X(_02738_));
 sky130_fd_sc_hd__inv_2 _17433_ (.A(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__buf_2 _17434_ (.A(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__buf_2 _17435_ (.A(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__a22oi_4 _17436_ (.A1(\CPU_Xreg_value_a4[23][0] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][0] ),
    .B2(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__or4_4 _17437_ (.A(_02662_),
    .B(_02658_),
    .C(_02676_),
    .D(_02653_),
    .X(_02743_));
 sky130_fd_sc_hd__buf_2 _17438_ (.A(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__buf_2 _17439_ (.A(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__or4_4 _17440_ (.A(_02662_),
    .B(_02702_),
    .C(_02676_),
    .D(_02678_),
    .X(_02746_));
 sky130_fd_sc_hd__buf_2 _17441_ (.A(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_2 _17442_ (.A(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__o22a_4 _17443_ (.A1(_08612_),
    .A2(_02745_),
    .B1(_07533_),
    .B2(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__and4_4 _17444_ (.A(_02726_),
    .B(_02733_),
    .C(_02742_),
    .D(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__or4_4 _17445_ (.A(_02664_),
    .B(_02658_),
    .C(_02690_),
    .D(_02677_),
    .X(_02751_));
 sky130_fd_sc_hd__buf_2 _17446_ (.A(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__buf_2 _17447_ (.A(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__or2_4 _17448_ (.A(_02663_),
    .B(_02657_),
    .X(_02754_));
 sky130_fd_sc_hd__or4_4 _17449_ (.A(_02650_),
    .B(_02646_),
    .C(_02754_),
    .D(_02678_),
    .X(_02755_));
 sky130_fd_sc_hd__buf_2 _17450_ (.A(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__buf_2 _17451_ (.A(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__o22a_4 _17452_ (.A1(_01654_),
    .A2(_02753_),
    .B1(_07733_),
    .B2(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__inv_2 _17453_ (.A(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__or4_4 _17454_ (.A(_02650_),
    .B(_02646_),
    .C(_02754_),
    .D(_02652_),
    .X(_02760_));
 sky130_fd_sc_hd__buf_2 _17455_ (.A(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__buf_2 _17456_ (.A(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__or4_4 _17457_ (.A(_02664_),
    .B(_02658_),
    .C(_02690_),
    .D(_02652_),
    .X(_02763_));
 sky130_fd_sc_hd__inv_2 _17458_ (.A(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__buf_2 _17459_ (.A(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__buf_2 _17460_ (.A(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__a2bb2o_4 _17461_ (.A1_N(_09130_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][0] ),
    .B2(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__or2_4 _17462_ (.A(_02663_),
    .B(_02695_),
    .X(_02768_));
 sky130_fd_sc_hd__or4_4 _17463_ (.A(_02650_),
    .B(_02646_),
    .C(_02768_),
    .D(_02677_),
    .X(_02769_));
 sky130_fd_sc_hd__inv_2 _17464_ (.A(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__buf_2 _17465_ (.A(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_2 _17466_ (.A(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__or4_4 _17467_ (.A(_02661_),
    .B(_02658_),
    .C(_02690_),
    .D(_02677_),
    .X(_02773_));
 sky130_fd_sc_hd__inv_2 _17468_ (.A(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__buf_2 _17469_ (.A(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__or2_4 _17470_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .B(_02657_),
    .X(_02776_));
 sky130_fd_sc_hd__or4_4 _17471_ (.A(_02649_),
    .B(_02645_),
    .C(_02776_),
    .D(_02652_),
    .X(_02777_));
 sky130_fd_sc_hd__buf_2 _17472_ (.A(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__buf_2 _17473_ (.A(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_2 _17474_ (.A(_02651_),
    .X(_02780_));
 sky130_fd_sc_hd__or4_4 _17475_ (.A(_02661_),
    .B(_02696_),
    .C(_02683_),
    .D(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__inv_2 _17476_ (.A(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__buf_2 _17477_ (.A(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__buf_2 _17478_ (.A(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__a2bb2o_4 _17479_ (.A1_N(_08445_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][0] ),
    .B2(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a211o_4 _17480_ (.A1(\CPU_Xreg_value_a4[13][0] ),
    .A2(_02772_),
    .B1(_02775_),
    .C1(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__inv_2 _17481_ (.A(\CPU_Xreg_value_a4[18][0] ),
    .Y(_02787_));
 sky130_fd_sc_hd__or4_4 _17482_ (.A(_02661_),
    .B(_02657_),
    .C(_02684_),
    .D(_02780_),
    .X(_02788_));
 sky130_fd_sc_hd__buf_2 _17483_ (.A(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__buf_2 _17484_ (.A(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__or4_4 _17485_ (.A(_02663_),
    .B(_02695_),
    .C(_02689_),
    .D(_02651_),
    .X(_02791_));
 sky130_fd_sc_hd__inv_2 _17486_ (.A(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__buf_2 _17487_ (.A(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__buf_2 _17488_ (.A(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__a2bb2o_4 _17489_ (.A1_N(_02787_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][0] ),
    .B2(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__or4_4 _17490_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .B(_02657_),
    .C(_02683_),
    .D(_02677_),
    .X(_02796_));
 sky130_fd_sc_hd__buf_2 _17491_ (.A(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__buf_2 _17492_ (.A(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__or4_4 _17493_ (.A(_02649_),
    .B(_02645_),
    .C(_02776_),
    .D(_02677_),
    .X(_02799_));
 sky130_fd_sc_hd__buf_2 _17494_ (.A(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__buf_2 _17495_ (.A(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__o22a_4 _17496_ (.A1(_01671_),
    .A2(_02798_),
    .B1(_06982_),
    .B2(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__inv_2 _17497_ (.A(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__or4_4 _17498_ (.A(_02649_),
    .B(_02645_),
    .C(_02706_),
    .D(_02780_),
    .X(_02804_));
 sky130_fd_sc_hd__buf_2 _17499_ (.A(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__buf_2 _17500_ (.A(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__or4_4 _17501_ (.A(\CPU_rf_rd_index2_a2[3] ),
    .B(_02696_),
    .C(_02689_),
    .D(_02780_),
    .X(_02807_));
 sky130_fd_sc_hd__inv_2 _17502_ (.A(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__buf_2 _17503_ (.A(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__buf_2 _17504_ (.A(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a2bb2o_4 _17505_ (.A1_N(_08804_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][0] ),
    .B2(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__or4_4 _17506_ (.A(_02663_),
    .B(_02657_),
    .C(_02675_),
    .D(_02780_),
    .X(_02812_));
 sky130_fd_sc_hd__buf_2 _17507_ (.A(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__buf_2 _17508_ (.A(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__or4_4 _17509_ (.A(_02649_),
    .B(_02645_),
    .C(_02768_),
    .D(_02780_),
    .X(_02815_));
 sky130_fd_sc_hd__inv_2 _17510_ (.A(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__buf_2 _17511_ (.A(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_2 _17512_ (.A(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__a2bb2o_4 _17513_ (.A1_N(_09322_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][0] ),
    .B2(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__or4_4 _17514_ (.A(_02795_),
    .B(_02803_),
    .C(_02811_),
    .D(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__or4_4 _17515_ (.A(_02759_),
    .B(_02767_),
    .C(_02786_),
    .D(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__inv_2 _17516_ (.A(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__buf_2 _17517_ (.A(_02775_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_2 _17518_ (.A(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__a32o_4 _17519_ (.A1(_02718_),
    .A2(_02750_),
    .A3(_02822_),
    .B1(_06142_),
    .B2(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__inv_2 _17520_ (.A(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o22a_4 _17521_ (.A1(_06979_),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02826_),
    .X(\CPU_src2_value_a2[0] ));
 sky130_fd_sc_hd__o22a_4 _17522_ (.A1(_07186_),
    .A2(_02682_),
    .B1(_07817_),
    .B2(_02687_),
    .X(_02827_));
 sky130_fd_sc_hd__a22oi_4 _17523_ (.A1(\CPU_Xreg_value_a4[16][1] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][1] ),
    .B2(_02700_),
    .Y(_02828_));
 sky130_fd_sc_hd__o22a_4 _17524_ (.A1(_07445_),
    .A2(_02705_),
    .B1(_01724_),
    .B2(_02709_),
    .X(_02829_));
 sky130_fd_sc_hd__o22a_4 _17525_ (.A1(_01734_),
    .A2(_02713_),
    .B1(_07900_),
    .B2(_02716_),
    .X(_02830_));
 sky130_fd_sc_hd__and4_4 _17526_ (.A(_02827_),
    .B(_02828_),
    .C(_02829_),
    .D(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__o22a_4 _17527_ (.A1(_09238_),
    .A2(_02722_),
    .B1(_01725_),
    .B2(_02725_),
    .X(_02832_));
 sky130_fd_sc_hd__o22a_4 _17528_ (.A1(_08268_),
    .A2(_02729_),
    .B1(_08182_),
    .B2(_02732_),
    .X(_02833_));
 sky130_fd_sc_hd__a22oi_4 _17529_ (.A1(\CPU_Xreg_value_a4[23][1] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][1] ),
    .B2(_02741_),
    .Y(_02834_));
 sky130_fd_sc_hd__o22a_4 _17530_ (.A1(_08610_),
    .A2(_02745_),
    .B1(_07531_),
    .B2(_02748_),
    .X(_02835_));
 sky130_fd_sc_hd__and4_4 _17531_ (.A(_02832_),
    .B(_02833_),
    .C(_02834_),
    .D(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__o22a_4 _17532_ (.A1(_01719_),
    .A2(_02753_),
    .B1(_01738_),
    .B2(_02757_),
    .X(_02837_));
 sky130_fd_sc_hd__inv_2 _17533_ (.A(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__inv_2 _17534_ (.A(\CPU_Xreg_value_a4[25][1] ),
    .Y(_02839_));
 sky130_fd_sc_hd__a2bb2o_4 _17535_ (.A1_N(_02839_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][1] ),
    .B2(_02766_),
    .X(_02840_));
 sky130_fd_sc_hd__inv_2 _17536_ (.A(\CPU_Xreg_value_a4[17][1] ),
    .Y(_02841_));
 sky130_fd_sc_hd__a2bb2o_4 _17537_ (.A1_N(_02841_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][1] ),
    .B2(_02784_),
    .X(_02842_));
 sky130_fd_sc_hd__a211o_4 _17538_ (.A1(\CPU_Xreg_value_a4[13][1] ),
    .A2(_02772_),
    .B1(_02775_),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a2bb2o_4 _17539_ (.A1_N(_08527_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][1] ),
    .B2(_02794_),
    .X(_02844_));
 sky130_fd_sc_hd__o22a_4 _17540_ (.A1(_07098_),
    .A2(_02798_),
    .B1(_01733_),
    .B2(_02801_),
    .X(_02845_));
 sky130_fd_sc_hd__inv_2 _17541_ (.A(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__inv_2 _17542_ (.A(\CPU_Xreg_value_a4[21][1] ),
    .Y(_02847_));
 sky130_fd_sc_hd__a2bb2o_4 _17543_ (.A1_N(_02847_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][1] ),
    .B2(_02810_),
    .X(_02848_));
 sky130_fd_sc_hd__a2bb2o_4 _17544_ (.A1_N(_09320_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][1] ),
    .B2(_02818_),
    .X(_02849_));
 sky130_fd_sc_hd__or4_4 _17545_ (.A(_02844_),
    .B(_02846_),
    .C(_02848_),
    .D(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__or4_4 _17546_ (.A(_02838_),
    .B(_02840_),
    .C(_02843_),
    .D(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__inv_2 _17547_ (.A(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__a32o_4 _17548_ (.A1(_02831_),
    .A2(_02836_),
    .A3(_02852_),
    .B1(_06141_),
    .B2(_02824_),
    .X(_02853_));
 sky130_fd_sc_hd__inv_2 _17549_ (.A(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__o22a_4 _17550_ (.A1(_06866_),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02854_),
    .X(\CPU_src2_value_a2[1] ));
 sky130_fd_sc_hd__o22a_4 _17551_ (.A1(_01749_),
    .A2(_02682_),
    .B1(_01757_),
    .B2(_02687_),
    .X(_02855_));
 sky130_fd_sc_hd__a22oi_4 _17552_ (.A1(\CPU_Xreg_value_a4[16][2] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][2] ),
    .B2(_02700_),
    .Y(_02856_));
 sky130_fd_sc_hd__o22a_4 _17553_ (.A1(_07443_),
    .A2(_02705_),
    .B1(_07359_),
    .B2(_02709_),
    .X(_02857_));
 sky130_fd_sc_hd__o22a_4 _17554_ (.A1(_07275_),
    .A2(_02713_),
    .B1(_01755_),
    .B2(_02716_),
    .X(_02858_));
 sky130_fd_sc_hd__and4_4 _17555_ (.A(_02855_),
    .B(_02856_),
    .C(_02857_),
    .D(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__inv_2 _17556_ (.A(\CPU_Xreg_value_a4[26][2] ),
    .Y(_02860_));
 sky130_fd_sc_hd__o22a_4 _17557_ (.A1(_02860_),
    .A2(_02722_),
    .B1(_07983_),
    .B2(_02725_),
    .X(_02861_));
 sky130_fd_sc_hd__o22a_4 _17558_ (.A1(_08266_),
    .A2(_02729_),
    .B1(_08179_),
    .B2(_02732_),
    .X(_02862_));
 sky130_fd_sc_hd__a22oi_4 _17559_ (.A1(\CPU_Xreg_value_a4[23][2] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][2] ),
    .B2(_02741_),
    .Y(_02863_));
 sky130_fd_sc_hd__inv_2 _17560_ (.A(\CPU_Xreg_value_a4[19][2] ),
    .Y(_02864_));
 sky130_fd_sc_hd__o22a_4 _17561_ (.A1(_02864_),
    .A2(_02745_),
    .B1(_07528_),
    .B2(_02748_),
    .X(_02865_));
 sky130_fd_sc_hd__and4_4 _17562_ (.A(_02861_),
    .B(_02862_),
    .C(_02863_),
    .D(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__o22a_4 _17563_ (.A1(_01743_),
    .A2(_02753_),
    .B1(_01759_),
    .B2(_02757_),
    .X(_02867_));
 sky130_fd_sc_hd__inv_2 _17564_ (.A(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__inv_2 _17565_ (.A(\CPU_Xreg_value_a4[25][2] ),
    .Y(_02869_));
 sky130_fd_sc_hd__a2bb2o_4 _17566_ (.A1_N(_02869_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][2] ),
    .B2(_02766_),
    .X(_02870_));
 sky130_fd_sc_hd__inv_2 _17567_ (.A(\CPU_Xreg_value_a4[17][2] ),
    .Y(_02871_));
 sky130_fd_sc_hd__a2bb2o_4 _17568_ (.A1_N(_02871_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][2] ),
    .B2(_02784_),
    .X(_02872_));
 sky130_fd_sc_hd__a211o_4 _17569_ (.A1(\CPU_Xreg_value_a4[13][2] ),
    .A2(_02772_),
    .B1(_02775_),
    .C1(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__inv_2 _17570_ (.A(\CPU_Xreg_value_a4[18][2] ),
    .Y(_02874_));
 sky130_fd_sc_hd__a2bb2o_4 _17571_ (.A1_N(_02874_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][2] ),
    .B2(_02794_),
    .X(_02875_));
 sky130_fd_sc_hd__o22a_4 _17572_ (.A1(_01747_),
    .A2(_02798_),
    .B1(_01753_),
    .B2(_02801_),
    .X(_02876_));
 sky130_fd_sc_hd__inv_2 _17573_ (.A(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__a2bb2o_4 _17574_ (.A1_N(_08800_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][2] ),
    .B2(_02810_),
    .X(_02878_));
 sky130_fd_sc_hd__inv_2 _17575_ (.A(\CPU_Xreg_value_a4[27][2] ),
    .Y(_02879_));
 sky130_fd_sc_hd__a2bb2o_4 _17576_ (.A1_N(_02879_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][2] ),
    .B2(_02818_),
    .X(_02880_));
 sky130_fd_sc_hd__or4_4 _17577_ (.A(_02875_),
    .B(_02877_),
    .C(_02878_),
    .D(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__or4_4 _17578_ (.A(_02868_),
    .B(_02870_),
    .C(_02873_),
    .D(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__inv_2 _17579_ (.A(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__a32o_4 _17580_ (.A1(_02859_),
    .A2(_02866_),
    .A3(_02883_),
    .B1(_06139_),
    .B2(_02824_),
    .X(_02884_));
 sky130_fd_sc_hd__inv_2 _17581_ (.A(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__o22a_4 _17582_ (.A1(\CPU_result_a3[2] ),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02885_),
    .X(\CPU_src2_value_a2[2] ));
 sky130_fd_sc_hd__o22a_4 _17583_ (.A1(_01770_),
    .A2(_02682_),
    .B1(_07812_),
    .B2(_02687_),
    .X(_02886_));
 sky130_fd_sc_hd__a22oi_4 _17584_ (.A1(\CPU_Xreg_value_a4[16][3] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][3] ),
    .B2(_02700_),
    .Y(_02887_));
 sky130_fd_sc_hd__o22a_4 _17585_ (.A1(_01777_),
    .A2(_02705_),
    .B1(_01765_),
    .B2(_02709_),
    .X(_02888_));
 sky130_fd_sc_hd__o22a_4 _17586_ (.A1(_01775_),
    .A2(_02713_),
    .B1(_07896_),
    .B2(_02716_),
    .X(_02889_));
 sky130_fd_sc_hd__and4_4 _17587_ (.A(_02886_),
    .B(_02887_),
    .C(_02888_),
    .D(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__o22a_4 _17588_ (.A1(_09234_),
    .A2(_02722_),
    .B1(_07981_),
    .B2(_02725_),
    .X(_02891_));
 sky130_fd_sc_hd__o22a_4 _17589_ (.A1(_08264_),
    .A2(_02729_),
    .B1(_08176_),
    .B2(_02732_),
    .X(_02892_));
 sky130_fd_sc_hd__a22oi_4 _17590_ (.A1(\CPU_Xreg_value_a4[23][3] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][3] ),
    .B2(_02741_),
    .Y(_02893_));
 sky130_fd_sc_hd__inv_2 _17591_ (.A(\CPU_Xreg_value_a4[19][3] ),
    .Y(_02894_));
 sky130_fd_sc_hd__o22a_4 _17592_ (.A1(_02894_),
    .A2(_02745_),
    .B1(_01780_),
    .B2(_02748_),
    .X(_02895_));
 sky130_fd_sc_hd__and4_4 _17593_ (.A(_02891_),
    .B(_02892_),
    .C(_02893_),
    .D(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__o22a_4 _17594_ (.A1(_07643_),
    .A2(_02753_),
    .B1(_07727_),
    .B2(_02757_),
    .X(_02897_));
 sky130_fd_sc_hd__inv_2 _17595_ (.A(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__a2bb2o_4 _17596_ (.A1_N(_09123_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][3] ),
    .B2(_02766_),
    .X(_02899_));
 sky130_fd_sc_hd__inv_2 _17597_ (.A(\CPU_Xreg_value_a4[17][3] ),
    .Y(_02900_));
 sky130_fd_sc_hd__a2bb2o_4 _17598_ (.A1_N(_02900_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][3] ),
    .B2(_02784_),
    .X(_02901_));
 sky130_fd_sc_hd__a211o_4 _17599_ (.A1(\CPU_Xreg_value_a4[13][3] ),
    .A2(_02772_),
    .B1(_02775_),
    .C1(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__inv_2 _17600_ (.A(\CPU_Xreg_value_a4[18][3] ),
    .Y(_02903_));
 sky130_fd_sc_hd__a2bb2o_4 _17601_ (.A1_N(_02903_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][3] ),
    .B2(_02794_),
    .X(_02904_));
 sky130_fd_sc_hd__o22a_4 _17602_ (.A1(_01768_),
    .A2(_02798_),
    .B1(_01774_),
    .B2(_02801_),
    .X(_02905_));
 sky130_fd_sc_hd__inv_2 _17603_ (.A(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__inv_2 _17604_ (.A(\CPU_Xreg_value_a4[21][3] ),
    .Y(_02907_));
 sky130_fd_sc_hd__a2bb2o_4 _17605_ (.A1_N(_02907_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][3] ),
    .B2(_02810_),
    .X(_02908_));
 sky130_fd_sc_hd__a2bb2o_4 _17606_ (.A1_N(_09316_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][3] ),
    .B2(_02818_),
    .X(_02909_));
 sky130_fd_sc_hd__or4_4 _17607_ (.A(_02904_),
    .B(_02906_),
    .C(_02908_),
    .D(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__or4_4 _17608_ (.A(_02898_),
    .B(_02899_),
    .C(_02902_),
    .D(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__inv_2 _17609_ (.A(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__a32o_4 _17610_ (.A1(_02890_),
    .A2(_02896_),
    .A3(_02912_),
    .B1(_06138_),
    .B2(_02824_),
    .X(_02913_));
 sky130_fd_sc_hd__inv_2 _17611_ (.A(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__o22a_4 _17612_ (.A1(\CPU_result_a3[3] ),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02914_),
    .X(\CPU_src2_value_a2[3] ));
 sky130_fd_sc_hd__o22a_4 _17613_ (.A1(_01794_),
    .A2(_02682_),
    .B1(_01805_),
    .B2(_02687_),
    .X(_02915_));
 sky130_fd_sc_hd__a22oi_4 _17614_ (.A1(\CPU_Xreg_value_a4[16][4] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][4] ),
    .B2(_02700_),
    .Y(_02916_));
 sky130_fd_sc_hd__o22a_4 _17615_ (.A1(_01801_),
    .A2(_02705_),
    .B1(_01787_),
    .B2(_02709_),
    .X(_02917_));
 sky130_fd_sc_hd__o22a_4 _17616_ (.A1(_01799_),
    .A2(_02713_),
    .B1(_01802_),
    .B2(_02716_),
    .X(_02918_));
 sky130_fd_sc_hd__and4_4 _17617_ (.A(_02915_),
    .B(_02916_),
    .C(_02917_),
    .D(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__o22a_4 _17618_ (.A1(_09231_),
    .A2(_02722_),
    .B1(_01788_),
    .B2(_02725_),
    .X(_02920_));
 sky130_fd_sc_hd__o22a_4 _17619_ (.A1(_01804_),
    .A2(_02729_),
    .B1(_01793_),
    .B2(_02732_),
    .X(_02921_));
 sky130_fd_sc_hd__a22oi_4 _17620_ (.A1(\CPU_Xreg_value_a4[23][4] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][4] ),
    .B2(_02741_),
    .Y(_02922_));
 sky130_fd_sc_hd__o22a_4 _17621_ (.A1(_08603_),
    .A2(_02745_),
    .B1(_01808_),
    .B2(_02748_),
    .X(_02923_));
 sky130_fd_sc_hd__and4_4 _17622_ (.A(_02920_),
    .B(_02921_),
    .C(_02922_),
    .D(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__o22a_4 _17623_ (.A1(_01785_),
    .A2(_02753_),
    .B1(_01807_),
    .B2(_02757_),
    .X(_02925_));
 sky130_fd_sc_hd__inv_2 _17624_ (.A(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__a2bb2o_4 _17625_ (.A1_N(_09121_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][4] ),
    .B2(_02766_),
    .X(_02927_));
 sky130_fd_sc_hd__buf_2 _17626_ (.A(_02774_),
    .X(_02928_));
 sky130_fd_sc_hd__buf_2 _17627_ (.A(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__a2bb2o_4 _17628_ (.A1_N(_08435_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][4] ),
    .B2(_02784_),
    .X(_02930_));
 sky130_fd_sc_hd__a211o_4 _17629_ (.A1(\CPU_Xreg_value_a4[13][4] ),
    .A2(_02772_),
    .B1(_02929_),
    .C1(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__a2bb2o_4 _17630_ (.A1_N(_08520_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][4] ),
    .B2(_02794_),
    .X(_02932_));
 sky130_fd_sc_hd__o22a_4 _17631_ (.A1(_01791_),
    .A2(_02798_),
    .B1(_01798_),
    .B2(_02801_),
    .X(_02933_));
 sky130_fd_sc_hd__inv_2 _17632_ (.A(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__a2bb2o_4 _17633_ (.A1_N(_08796_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][4] ),
    .B2(_02810_),
    .X(_02935_));
 sky130_fd_sc_hd__a2bb2o_4 _17634_ (.A1_N(_09314_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][4] ),
    .B2(_02818_),
    .X(_02936_));
 sky130_fd_sc_hd__or4_4 _17635_ (.A(_02932_),
    .B(_02934_),
    .C(_02935_),
    .D(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__or4_4 _17636_ (.A(_02926_),
    .B(_02927_),
    .C(_02931_),
    .D(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__inv_2 _17637_ (.A(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__a32o_4 _17638_ (.A1(_02919_),
    .A2(_02924_),
    .A3(_02939_),
    .B1(_06137_),
    .B2(_02824_),
    .X(_02940_));
 sky130_fd_sc_hd__inv_2 _17639_ (.A(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__o22a_4 _17640_ (.A1(\CPU_result_a3[4] ),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02941_),
    .X(\CPU_src2_value_a2[4] ));
 sky130_fd_sc_hd__o22a_4 _17641_ (.A1(_01823_),
    .A2(_02682_),
    .B1(_01834_),
    .B2(_02687_),
    .X(_02942_));
 sky130_fd_sc_hd__a22oi_4 _17642_ (.A1(\CPU_Xreg_value_a4[16][5] ),
    .A2(_02694_),
    .B1(\CPU_Xreg_value_a4[30][5] ),
    .B2(_02700_),
    .Y(_02943_));
 sky130_fd_sc_hd__o22a_4 _17643_ (.A1(_01830_),
    .A2(_02705_),
    .B1(_01815_),
    .B2(_02709_),
    .X(_02944_));
 sky130_fd_sc_hd__o22a_4 _17644_ (.A1(_01828_),
    .A2(_02713_),
    .B1(_01831_),
    .B2(_02716_),
    .X(_02945_));
 sky130_fd_sc_hd__and4_4 _17645_ (.A(_02942_),
    .B(_02943_),
    .C(_02944_),
    .D(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__inv_2 _17646_ (.A(\CPU_Xreg_value_a4[26][5] ),
    .Y(_02947_));
 sky130_fd_sc_hd__o22a_4 _17647_ (.A1(_02947_),
    .A2(_02722_),
    .B1(_01816_),
    .B2(_02725_),
    .X(_02948_));
 sky130_fd_sc_hd__o22a_4 _17648_ (.A1(_01833_),
    .A2(_02729_),
    .B1(_01822_),
    .B2(_02732_),
    .X(_02949_));
 sky130_fd_sc_hd__a22oi_4 _17649_ (.A1(\CPU_Xreg_value_a4[23][5] ),
    .A2(_02737_),
    .B1(\CPU_Xreg_value_a4[31][5] ),
    .B2(_02741_),
    .Y(_02950_));
 sky130_fd_sc_hd__inv_2 _17650_ (.A(\CPU_Xreg_value_a4[19][5] ),
    .Y(_02951_));
 sky130_fd_sc_hd__o22a_4 _17651_ (.A1(_02951_),
    .A2(_02745_),
    .B1(_01837_),
    .B2(_02748_),
    .X(_02952_));
 sky130_fd_sc_hd__and4_4 _17652_ (.A(_02948_),
    .B(_02949_),
    .C(_02950_),
    .D(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o22a_4 _17653_ (.A1(_01813_),
    .A2(_02753_),
    .B1(_01836_),
    .B2(_02757_),
    .X(_02954_));
 sky130_fd_sc_hd__inv_2 _17654_ (.A(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__inv_2 _17655_ (.A(\CPU_Xreg_value_a4[25][5] ),
    .Y(_02956_));
 sky130_fd_sc_hd__a2bb2o_4 _17656_ (.A1_N(_02956_),
    .A2_N(_02762_),
    .B1(\CPU_Xreg_value_a4[24][5] ),
    .B2(_02766_),
    .X(_02957_));
 sky130_fd_sc_hd__inv_2 _17657_ (.A(\CPU_Xreg_value_a4[17][5] ),
    .Y(_02958_));
 sky130_fd_sc_hd__a2bb2o_4 _17658_ (.A1_N(_02958_),
    .A2_N(_02779_),
    .B1(\CPU_Xreg_value_a4[22][5] ),
    .B2(_02784_),
    .X(_02959_));
 sky130_fd_sc_hd__a211o_4 _17659_ (.A1(\CPU_Xreg_value_a4[13][5] ),
    .A2(_02772_),
    .B1(_02929_),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__inv_2 _17660_ (.A(\CPU_Xreg_value_a4[18][5] ),
    .Y(_02961_));
 sky130_fd_sc_hd__a2bb2o_4 _17661_ (.A1_N(_02961_),
    .A2_N(_02790_),
    .B1(\CPU_Xreg_value_a4[28][5] ),
    .B2(_02794_),
    .X(_02962_));
 sky130_fd_sc_hd__o22a_4 _17662_ (.A1(_01819_),
    .A2(_02798_),
    .B1(_01827_),
    .B2(_02801_),
    .X(_02963_));
 sky130_fd_sc_hd__inv_2 _17663_ (.A(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__inv_2 _17664_ (.A(\CPU_Xreg_value_a4[21][5] ),
    .Y(_02965_));
 sky130_fd_sc_hd__a2bb2o_4 _17665_ (.A1_N(_02965_),
    .A2_N(_02806_),
    .B1(\CPU_Xreg_value_a4[20][5] ),
    .B2(_02810_),
    .X(_02966_));
 sky130_fd_sc_hd__inv_2 _17666_ (.A(\CPU_Xreg_value_a4[27][5] ),
    .Y(_02967_));
 sky130_fd_sc_hd__a2bb2o_4 _17667_ (.A1_N(_02967_),
    .A2_N(_02814_),
    .B1(\CPU_Xreg_value_a4[29][5] ),
    .B2(_02818_),
    .X(_02968_));
 sky130_fd_sc_hd__or4_4 _17668_ (.A(_02962_),
    .B(_02964_),
    .C(_02966_),
    .D(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__or4_4 _17669_ (.A(_02955_),
    .B(_02957_),
    .C(_02960_),
    .D(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__inv_2 _17670_ (.A(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__a32o_4 _17671_ (.A1(_02946_),
    .A2(_02953_),
    .A3(_02971_),
    .B1(_06136_),
    .B2(_02824_),
    .X(_02972_));
 sky130_fd_sc_hd__inv_2 _17672_ (.A(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__o22a_4 _17673_ (.A1(\CPU_result_a3[5] ),
    .A2(_02670_),
    .B1(_02673_),
    .B2(_02973_),
    .X(\CPU_src2_value_a2[5] ));
 sky130_fd_sc_hd__buf_2 _17674_ (.A(_02669_),
    .X(_02974_));
 sky130_fd_sc_hd__buf_2 _17675_ (.A(_02672_),
    .X(_02975_));
 sky130_fd_sc_hd__buf_2 _17676_ (.A(_02681_),
    .X(_02976_));
 sky130_fd_sc_hd__buf_2 _17677_ (.A(_02686_),
    .X(_02977_));
 sky130_fd_sc_hd__o22a_4 _17678_ (.A1(_01856_),
    .A2(_02976_),
    .B1(_01873_),
    .B2(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_2 _17679_ (.A(_02693_),
    .X(_02979_));
 sky130_fd_sc_hd__buf_2 _17680_ (.A(_02699_),
    .X(_02980_));
 sky130_fd_sc_hd__a22oi_4 _17681_ (.A1(\CPU_Xreg_value_a4[16][6] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][6] ),
    .B2(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__buf_2 _17682_ (.A(_02704_),
    .X(_02982_));
 sky130_fd_sc_hd__buf_2 _17683_ (.A(_02708_),
    .X(_02983_));
 sky130_fd_sc_hd__o22a_4 _17684_ (.A1(_01866_),
    .A2(_02982_),
    .B1(_01846_),
    .B2(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__buf_2 _17685_ (.A(_02712_),
    .X(_02985_));
 sky130_fd_sc_hd__buf_2 _17686_ (.A(_02715_),
    .X(_02986_));
 sky130_fd_sc_hd__o22a_4 _17687_ (.A1(_01863_),
    .A2(_02985_),
    .B1(_01868_),
    .B2(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__and4_4 _17688_ (.A(_02978_),
    .B(_02981_),
    .C(_02984_),
    .D(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__inv_2 _17689_ (.A(\CPU_Xreg_value_a4[26][6] ),
    .Y(_02989_));
 sky130_fd_sc_hd__buf_2 _17690_ (.A(_02721_),
    .X(_02990_));
 sky130_fd_sc_hd__buf_2 _17691_ (.A(_02724_),
    .X(_02991_));
 sky130_fd_sc_hd__o22a_4 _17692_ (.A1(_02989_),
    .A2(_02990_),
    .B1(_01848_),
    .B2(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__buf_2 _17693_ (.A(_02728_),
    .X(_02993_));
 sky130_fd_sc_hd__buf_2 _17694_ (.A(_02731_),
    .X(_02994_));
 sky130_fd_sc_hd__o22a_4 _17695_ (.A1(_01871_),
    .A2(_02993_),
    .B1(_01854_),
    .B2(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__buf_2 _17696_ (.A(_02736_),
    .X(_02996_));
 sky130_fd_sc_hd__buf_2 _17697_ (.A(_02740_),
    .X(_02997_));
 sky130_fd_sc_hd__a22oi_4 _17698_ (.A1(\CPU_Xreg_value_a4[23][6] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][6] ),
    .B2(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__inv_2 _17699_ (.A(\CPU_Xreg_value_a4[19][6] ),
    .Y(_02999_));
 sky130_fd_sc_hd__buf_2 _17700_ (.A(_02744_),
    .X(_03000_));
 sky130_fd_sc_hd__buf_2 _17701_ (.A(_02747_),
    .X(_03001_));
 sky130_fd_sc_hd__o22a_4 _17702_ (.A1(_02999_),
    .A2(_03000_),
    .B1(_01878_),
    .B2(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__and4_4 _17703_ (.A(_02992_),
    .B(_02995_),
    .C(_02998_),
    .D(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__buf_2 _17704_ (.A(_02752_),
    .X(_03004_));
 sky130_fd_sc_hd__buf_2 _17705_ (.A(_02756_),
    .X(_03005_));
 sky130_fd_sc_hd__o22a_4 _17706_ (.A1(_01844_),
    .A2(_03004_),
    .B1(_01876_),
    .B2(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__inv_2 _17707_ (.A(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__inv_2 _17708_ (.A(\CPU_Xreg_value_a4[25][6] ),
    .Y(_03008_));
 sky130_fd_sc_hd__buf_2 _17709_ (.A(_02761_),
    .X(_03009_));
 sky130_fd_sc_hd__buf_2 _17710_ (.A(_02765_),
    .X(_03010_));
 sky130_fd_sc_hd__a2bb2o_4 _17711_ (.A1_N(_03008_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][6] ),
    .B2(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_2 _17712_ (.A(_02771_),
    .X(_03012_));
 sky130_fd_sc_hd__inv_2 _17713_ (.A(\CPU_Xreg_value_a4[17][6] ),
    .Y(_03013_));
 sky130_fd_sc_hd__buf_2 _17714_ (.A(_02778_),
    .X(_03014_));
 sky130_fd_sc_hd__buf_2 _17715_ (.A(_02783_),
    .X(_03015_));
 sky130_fd_sc_hd__a2bb2o_4 _17716_ (.A1_N(_03013_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][6] ),
    .B2(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__a211o_4 _17717_ (.A1(\CPU_Xreg_value_a4[13][6] ),
    .A2(_03012_),
    .B1(_02929_),
    .C1(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__inv_2 _17718_ (.A(\CPU_Xreg_value_a4[18][6] ),
    .Y(_03018_));
 sky130_fd_sc_hd__buf_2 _17719_ (.A(_02789_),
    .X(_03019_));
 sky130_fd_sc_hd__buf_2 _17720_ (.A(_02793_),
    .X(_03020_));
 sky130_fd_sc_hd__a2bb2o_4 _17721_ (.A1_N(_03018_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][6] ),
    .B2(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__buf_2 _17722_ (.A(_02797_),
    .X(_03022_));
 sky130_fd_sc_hd__buf_2 _17723_ (.A(_02800_),
    .X(_03023_));
 sky130_fd_sc_hd__o22a_4 _17724_ (.A1(_01852_),
    .A2(_03022_),
    .B1(_01861_),
    .B2(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__inv_2 _17725_ (.A(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__inv_2 _17726_ (.A(\CPU_Xreg_value_a4[21][6] ),
    .Y(_03026_));
 sky130_fd_sc_hd__buf_2 _17727_ (.A(_02805_),
    .X(_03027_));
 sky130_fd_sc_hd__buf_2 _17728_ (.A(_02809_),
    .X(_03028_));
 sky130_fd_sc_hd__a2bb2o_4 _17729_ (.A1_N(_03026_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][6] ),
    .B2(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__inv_2 _17730_ (.A(\CPU_Xreg_value_a4[27][6] ),
    .Y(_03030_));
 sky130_fd_sc_hd__buf_2 _17731_ (.A(_02813_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_2 _17732_ (.A(_02817_),
    .X(_03032_));
 sky130_fd_sc_hd__a2bb2o_4 _17733_ (.A1_N(_03030_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][6] ),
    .B2(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__or4_4 _17734_ (.A(_03021_),
    .B(_03025_),
    .C(_03029_),
    .D(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__or4_4 _17735_ (.A(_03007_),
    .B(_03011_),
    .C(_03017_),
    .D(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__inv_2 _17736_ (.A(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__buf_2 _17737_ (.A(_02823_),
    .X(_03037_));
 sky130_fd_sc_hd__a32o_4 _17738_ (.A1(_02988_),
    .A2(_03003_),
    .A3(_03036_),
    .B1(_06135_),
    .B2(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__inv_2 _17739_ (.A(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__o22a_4 _17740_ (.A1(_06826_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03039_),
    .X(\CPU_src2_value_a2[6] ));
 sky130_fd_sc_hd__o22a_4 _17741_ (.A1(_01897_),
    .A2(_02976_),
    .B1(_01908_),
    .B2(_02977_),
    .X(_03040_));
 sky130_fd_sc_hd__a22oi_4 _17742_ (.A1(\CPU_Xreg_value_a4[16][7] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][7] ),
    .B2(_02980_),
    .Y(_03041_));
 sky130_fd_sc_hd__o22a_4 _17743_ (.A1(_01904_),
    .A2(_02982_),
    .B1(_01889_),
    .B2(_02983_),
    .X(_03042_));
 sky130_fd_sc_hd__o22a_4 _17744_ (.A1(_01902_),
    .A2(_02985_),
    .B1(_01905_),
    .B2(_02986_),
    .X(_03043_));
 sky130_fd_sc_hd__and4_4 _17745_ (.A(_03040_),
    .B(_03041_),
    .C(_03042_),
    .D(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__inv_2 _17746_ (.A(\CPU_Xreg_value_a4[26][7] ),
    .Y(_03045_));
 sky130_fd_sc_hd__o22a_4 _17747_ (.A1(_03045_),
    .A2(_02990_),
    .B1(_01890_),
    .B2(_02991_),
    .X(_03046_));
 sky130_fd_sc_hd__o22a_4 _17748_ (.A1(_01907_),
    .A2(_02993_),
    .B1(_01896_),
    .B2(_02994_),
    .X(_03047_));
 sky130_fd_sc_hd__a22oi_4 _17749_ (.A1(\CPU_Xreg_value_a4[23][7] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][7] ),
    .B2(_02997_),
    .Y(_03048_));
 sky130_fd_sc_hd__inv_2 _17750_ (.A(\CPU_Xreg_value_a4[19][7] ),
    .Y(_03049_));
 sky130_fd_sc_hd__o22a_4 _17751_ (.A1(_03049_),
    .A2(_03000_),
    .B1(_01911_),
    .B2(_03001_),
    .X(_03050_));
 sky130_fd_sc_hd__and4_4 _17752_ (.A(_03046_),
    .B(_03047_),
    .C(_03048_),
    .D(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__o22a_4 _17753_ (.A1(_01885_),
    .A2(_03004_),
    .B1(_01910_),
    .B2(_03005_),
    .X(_03052_));
 sky130_fd_sc_hd__inv_2 _17754_ (.A(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__inv_2 _17755_ (.A(\CPU_Xreg_value_a4[25][7] ),
    .Y(_03054_));
 sky130_fd_sc_hd__a2bb2o_4 _17756_ (.A1_N(_03054_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][7] ),
    .B2(_03010_),
    .X(_03055_));
 sky130_fd_sc_hd__inv_2 _17757_ (.A(\CPU_Xreg_value_a4[17][7] ),
    .Y(_03056_));
 sky130_fd_sc_hd__a2bb2o_4 _17758_ (.A1_N(_03056_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][7] ),
    .B2(_03015_),
    .X(_03057_));
 sky130_fd_sc_hd__a211o_4 _17759_ (.A1(\CPU_Xreg_value_a4[13][7] ),
    .A2(_03012_),
    .B1(_02929_),
    .C1(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__inv_2 _17760_ (.A(\CPU_Xreg_value_a4[18][7] ),
    .Y(_03059_));
 sky130_fd_sc_hd__a2bb2o_4 _17761_ (.A1_N(_03059_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][7] ),
    .B2(_03020_),
    .X(_03060_));
 sky130_fd_sc_hd__o22a_4 _17762_ (.A1(_01893_),
    .A2(_03022_),
    .B1(_01901_),
    .B2(_03023_),
    .X(_03061_));
 sky130_fd_sc_hd__inv_2 _17763_ (.A(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__inv_2 _17764_ (.A(\CPU_Xreg_value_a4[21][7] ),
    .Y(_03063_));
 sky130_fd_sc_hd__a2bb2o_4 _17765_ (.A1_N(_03063_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][7] ),
    .B2(_03028_),
    .X(_03064_));
 sky130_fd_sc_hd__inv_2 _17766_ (.A(\CPU_Xreg_value_a4[27][7] ),
    .Y(_03065_));
 sky130_fd_sc_hd__a2bb2o_4 _17767_ (.A1_N(_03065_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][7] ),
    .B2(_03032_),
    .X(_03066_));
 sky130_fd_sc_hd__or4_4 _17768_ (.A(_03060_),
    .B(_03062_),
    .C(_03064_),
    .D(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__or4_4 _17769_ (.A(_03053_),
    .B(_03055_),
    .C(_03058_),
    .D(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__inv_2 _17770_ (.A(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__a32o_4 _17771_ (.A1(_03044_),
    .A2(_03051_),
    .A3(_03069_),
    .B1(_06134_),
    .B2(_03037_),
    .X(_03070_));
 sky130_fd_sc_hd__inv_2 _17772_ (.A(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__o22a_4 _17773_ (.A1(_06818_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03071_),
    .X(\CPU_src2_value_a2[7] ));
 sky130_fd_sc_hd__o22a_4 _17774_ (.A1(_01925_),
    .A2(_02976_),
    .B1(_01936_),
    .B2(_02977_),
    .X(_03072_));
 sky130_fd_sc_hd__a22oi_4 _17775_ (.A1(\CPU_Xreg_value_a4[16][8] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][8] ),
    .B2(_02980_),
    .Y(_03073_));
 sky130_fd_sc_hd__o22a_4 _17776_ (.A1(_01932_),
    .A2(_02982_),
    .B1(_01918_),
    .B2(_02983_),
    .X(_03074_));
 sky130_fd_sc_hd__o22a_4 _17777_ (.A1(_01930_),
    .A2(_02985_),
    .B1(_01933_),
    .B2(_02986_),
    .X(_03075_));
 sky130_fd_sc_hd__and4_4 _17778_ (.A(_03072_),
    .B(_03073_),
    .C(_03074_),
    .D(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__inv_2 _17779_ (.A(\CPU_Xreg_value_a4[26][8] ),
    .Y(_03077_));
 sky130_fd_sc_hd__o22a_4 _17780_ (.A1(_03077_),
    .A2(_02990_),
    .B1(_01919_),
    .B2(_02991_),
    .X(_03078_));
 sky130_fd_sc_hd__o22a_4 _17781_ (.A1(_01935_),
    .A2(_02993_),
    .B1(_01924_),
    .B2(_02994_),
    .X(_03079_));
 sky130_fd_sc_hd__a22oi_4 _17782_ (.A1(\CPU_Xreg_value_a4[23][8] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][8] ),
    .B2(_02997_),
    .Y(_03080_));
 sky130_fd_sc_hd__inv_2 _17783_ (.A(\CPU_Xreg_value_a4[19][8] ),
    .Y(_03081_));
 sky130_fd_sc_hd__o22a_4 _17784_ (.A1(_03081_),
    .A2(_03000_),
    .B1(_01939_),
    .B2(_03001_),
    .X(_03082_));
 sky130_fd_sc_hd__and4_4 _17785_ (.A(_03078_),
    .B(_03079_),
    .C(_03080_),
    .D(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__o22a_4 _17786_ (.A1(_01916_),
    .A2(_03004_),
    .B1(_01938_),
    .B2(_03005_),
    .X(_03084_));
 sky130_fd_sc_hd__inv_2 _17787_ (.A(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__inv_2 _17788_ (.A(\CPU_Xreg_value_a4[25][8] ),
    .Y(_03086_));
 sky130_fd_sc_hd__a2bb2o_4 _17789_ (.A1_N(_03086_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][8] ),
    .B2(_03010_),
    .X(_03087_));
 sky130_fd_sc_hd__inv_2 _17790_ (.A(\CPU_Xreg_value_a4[17][8] ),
    .Y(_03088_));
 sky130_fd_sc_hd__a2bb2o_4 _17791_ (.A1_N(_03088_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][8] ),
    .B2(_03015_),
    .X(_03089_));
 sky130_fd_sc_hd__a211o_4 _17792_ (.A1(\CPU_Xreg_value_a4[13][8] ),
    .A2(_03012_),
    .B1(_02929_),
    .C1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__inv_2 _17793_ (.A(\CPU_Xreg_value_a4[18][8] ),
    .Y(_03091_));
 sky130_fd_sc_hd__a2bb2o_4 _17794_ (.A1_N(_03091_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][8] ),
    .B2(_03020_),
    .X(_03092_));
 sky130_fd_sc_hd__o22a_4 _17795_ (.A1(_01922_),
    .A2(_03022_),
    .B1(_01929_),
    .B2(_03023_),
    .X(_03093_));
 sky130_fd_sc_hd__inv_2 _17796_ (.A(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__inv_2 _17797_ (.A(\CPU_Xreg_value_a4[21][8] ),
    .Y(_03095_));
 sky130_fd_sc_hd__a2bb2o_4 _17798_ (.A1_N(_03095_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][8] ),
    .B2(_03028_),
    .X(_03096_));
 sky130_fd_sc_hd__inv_2 _17799_ (.A(\CPU_Xreg_value_a4[27][8] ),
    .Y(_03097_));
 sky130_fd_sc_hd__a2bb2o_4 _17800_ (.A1_N(_03097_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][8] ),
    .B2(_03032_),
    .X(_03098_));
 sky130_fd_sc_hd__or4_4 _17801_ (.A(_03092_),
    .B(_03094_),
    .C(_03096_),
    .D(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__or4_4 _17802_ (.A(_03085_),
    .B(_03087_),
    .C(_03090_),
    .D(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__inv_2 _17803_ (.A(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__a32o_4 _17804_ (.A1(_03076_),
    .A2(_03083_),
    .A3(_03101_),
    .B1(_06132_),
    .B2(_03037_),
    .X(_03102_));
 sky130_fd_sc_hd__inv_2 _17805_ (.A(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__o22a_4 _17806_ (.A1(_06797_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03103_),
    .X(\CPU_src2_value_a2[8] ));
 sky130_fd_sc_hd__o22a_4 _17807_ (.A1(_01953_),
    .A2(_02976_),
    .B1(_01964_),
    .B2(_02977_),
    .X(_03104_));
 sky130_fd_sc_hd__a22oi_4 _17808_ (.A1(\CPU_Xreg_value_a4[16][9] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][9] ),
    .B2(_02980_),
    .Y(_03105_));
 sky130_fd_sc_hd__o22a_4 _17809_ (.A1(_01960_),
    .A2(_02982_),
    .B1(_01946_),
    .B2(_02983_),
    .X(_03106_));
 sky130_fd_sc_hd__o22a_4 _17810_ (.A1(_01958_),
    .A2(_02985_),
    .B1(_01961_),
    .B2(_02986_),
    .X(_03107_));
 sky130_fd_sc_hd__and4_4 _17811_ (.A(_03104_),
    .B(_03105_),
    .C(_03106_),
    .D(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__inv_2 _17812_ (.A(\CPU_Xreg_value_a4[26][9] ),
    .Y(_03109_));
 sky130_fd_sc_hd__o22a_4 _17813_ (.A1(_03109_),
    .A2(_02990_),
    .B1(_01947_),
    .B2(_02991_),
    .X(_03110_));
 sky130_fd_sc_hd__o22a_4 _17814_ (.A1(_01963_),
    .A2(_02993_),
    .B1(_01952_),
    .B2(_02994_),
    .X(_03111_));
 sky130_fd_sc_hd__a22oi_4 _17815_ (.A1(\CPU_Xreg_value_a4[23][9] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][9] ),
    .B2(_02997_),
    .Y(_03112_));
 sky130_fd_sc_hd__inv_2 _17816_ (.A(\CPU_Xreg_value_a4[19][9] ),
    .Y(_03113_));
 sky130_fd_sc_hd__o22a_4 _17817_ (.A1(_03113_),
    .A2(_03000_),
    .B1(_01967_),
    .B2(_03001_),
    .X(_03114_));
 sky130_fd_sc_hd__and4_4 _17818_ (.A(_03110_),
    .B(_03111_),
    .C(_03112_),
    .D(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__o22a_4 _17819_ (.A1(_01944_),
    .A2(_03004_),
    .B1(_01966_),
    .B2(_03005_),
    .X(_03116_));
 sky130_fd_sc_hd__inv_2 _17820_ (.A(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__inv_2 _17821_ (.A(\CPU_Xreg_value_a4[25][9] ),
    .Y(_03118_));
 sky130_fd_sc_hd__a2bb2o_4 _17822_ (.A1_N(_03118_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][9] ),
    .B2(_03010_),
    .X(_03119_));
 sky130_fd_sc_hd__inv_2 _17823_ (.A(\CPU_Xreg_value_a4[17][9] ),
    .Y(_03120_));
 sky130_fd_sc_hd__a2bb2o_4 _17824_ (.A1_N(_03120_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][9] ),
    .B2(_03015_),
    .X(_03121_));
 sky130_fd_sc_hd__a211o_4 _17825_ (.A1(\CPU_Xreg_value_a4[13][9] ),
    .A2(_03012_),
    .B1(_02929_),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__inv_2 _17826_ (.A(\CPU_Xreg_value_a4[18][9] ),
    .Y(_03123_));
 sky130_fd_sc_hd__a2bb2o_4 _17827_ (.A1_N(_03123_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][9] ),
    .B2(_03020_),
    .X(_03124_));
 sky130_fd_sc_hd__o22a_4 _17828_ (.A1(_01950_),
    .A2(_03022_),
    .B1(_01957_),
    .B2(_03023_),
    .X(_03125_));
 sky130_fd_sc_hd__inv_2 _17829_ (.A(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__inv_2 _17830_ (.A(\CPU_Xreg_value_a4[21][9] ),
    .Y(_03127_));
 sky130_fd_sc_hd__a2bb2o_4 _17831_ (.A1_N(_03127_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][9] ),
    .B2(_03028_),
    .X(_03128_));
 sky130_fd_sc_hd__inv_2 _17832_ (.A(\CPU_Xreg_value_a4[27][9] ),
    .Y(_03129_));
 sky130_fd_sc_hd__a2bb2o_4 _17833_ (.A1_N(_03129_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][9] ),
    .B2(_03032_),
    .X(_03130_));
 sky130_fd_sc_hd__or4_4 _17834_ (.A(_03124_),
    .B(_03126_),
    .C(_03128_),
    .D(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__or4_4 _17835_ (.A(_03117_),
    .B(_03119_),
    .C(_03122_),
    .D(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__inv_2 _17836_ (.A(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__a32o_4 _17837_ (.A1(_03108_),
    .A2(_03115_),
    .A3(_03133_),
    .B1(_06131_),
    .B2(_03037_),
    .X(_03134_));
 sky130_fd_sc_hd__inv_2 _17838_ (.A(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__o22a_4 _17839_ (.A1(_06789_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03135_),
    .X(\CPU_src2_value_a2[9] ));
 sky130_fd_sc_hd__o22a_4 _17840_ (.A1(_01981_),
    .A2(_02976_),
    .B1(_01992_),
    .B2(_02977_),
    .X(_03136_));
 sky130_fd_sc_hd__a22oi_4 _17841_ (.A1(\CPU_Xreg_value_a4[16][10] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][10] ),
    .B2(_02980_),
    .Y(_03137_));
 sky130_fd_sc_hd__o22a_4 _17842_ (.A1(_01988_),
    .A2(_02982_),
    .B1(_01974_),
    .B2(_02983_),
    .X(_03138_));
 sky130_fd_sc_hd__o22a_4 _17843_ (.A1(_01986_),
    .A2(_02985_),
    .B1(_01989_),
    .B2(_02986_),
    .X(_03139_));
 sky130_fd_sc_hd__and4_4 _17844_ (.A(_03136_),
    .B(_03137_),
    .C(_03138_),
    .D(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__inv_2 _17845_ (.A(\CPU_Xreg_value_a4[26][10] ),
    .Y(_03141_));
 sky130_fd_sc_hd__o22a_4 _17846_ (.A1(_03141_),
    .A2(_02990_),
    .B1(_01975_),
    .B2(_02991_),
    .X(_03142_));
 sky130_fd_sc_hd__o22a_4 _17847_ (.A1(_01991_),
    .A2(_02993_),
    .B1(_01980_),
    .B2(_02994_),
    .X(_03143_));
 sky130_fd_sc_hd__a22oi_4 _17848_ (.A1(\CPU_Xreg_value_a4[23][10] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][10] ),
    .B2(_02997_),
    .Y(_03144_));
 sky130_fd_sc_hd__inv_2 _17849_ (.A(\CPU_Xreg_value_a4[19][10] ),
    .Y(_03145_));
 sky130_fd_sc_hd__o22a_4 _17850_ (.A1(_03145_),
    .A2(_03000_),
    .B1(_01995_),
    .B2(_03001_),
    .X(_03146_));
 sky130_fd_sc_hd__and4_4 _17851_ (.A(_03142_),
    .B(_03143_),
    .C(_03144_),
    .D(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__o22a_4 _17852_ (.A1(_01972_),
    .A2(_03004_),
    .B1(_01994_),
    .B2(_03005_),
    .X(_03148_));
 sky130_fd_sc_hd__inv_2 _17853_ (.A(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__inv_2 _17854_ (.A(\CPU_Xreg_value_a4[25][10] ),
    .Y(_03150_));
 sky130_fd_sc_hd__a2bb2o_4 _17855_ (.A1_N(_03150_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][10] ),
    .B2(_03010_),
    .X(_03151_));
 sky130_fd_sc_hd__buf_2 _17856_ (.A(_02928_),
    .X(_03152_));
 sky130_fd_sc_hd__inv_2 _17857_ (.A(\CPU_Xreg_value_a4[17][10] ),
    .Y(_03153_));
 sky130_fd_sc_hd__a2bb2o_4 _17858_ (.A1_N(_03153_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][10] ),
    .B2(_03015_),
    .X(_03154_));
 sky130_fd_sc_hd__a211o_4 _17859_ (.A1(\CPU_Xreg_value_a4[13][10] ),
    .A2(_03012_),
    .B1(_03152_),
    .C1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__inv_2 _17860_ (.A(\CPU_Xreg_value_a4[18][10] ),
    .Y(_03156_));
 sky130_fd_sc_hd__a2bb2o_4 _17861_ (.A1_N(_03156_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][10] ),
    .B2(_03020_),
    .X(_03157_));
 sky130_fd_sc_hd__o22a_4 _17862_ (.A1(_01978_),
    .A2(_03022_),
    .B1(_01985_),
    .B2(_03023_),
    .X(_03158_));
 sky130_fd_sc_hd__inv_2 _17863_ (.A(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__inv_2 _17864_ (.A(\CPU_Xreg_value_a4[21][10] ),
    .Y(_03160_));
 sky130_fd_sc_hd__a2bb2o_4 _17865_ (.A1_N(_03160_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][10] ),
    .B2(_03028_),
    .X(_03161_));
 sky130_fd_sc_hd__inv_2 _17866_ (.A(\CPU_Xreg_value_a4[27][10] ),
    .Y(_03162_));
 sky130_fd_sc_hd__a2bb2o_4 _17867_ (.A1_N(_03162_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][10] ),
    .B2(_03032_),
    .X(_03163_));
 sky130_fd_sc_hd__or4_4 _17868_ (.A(_03157_),
    .B(_03159_),
    .C(_03161_),
    .D(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__or4_4 _17869_ (.A(_03149_),
    .B(_03151_),
    .C(_03155_),
    .D(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__inv_2 _17870_ (.A(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a32o_4 _17871_ (.A1(_03140_),
    .A2(_03147_),
    .A3(_03166_),
    .B1(_06130_),
    .B2(_03037_),
    .X(_03167_));
 sky130_fd_sc_hd__inv_2 _17872_ (.A(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__o22a_4 _17873_ (.A1(_06776_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03168_),
    .X(\CPU_src2_value_a2[10] ));
 sky130_fd_sc_hd__o22a_4 _17874_ (.A1(_02010_),
    .A2(_02976_),
    .B1(_02021_),
    .B2(_02977_),
    .X(_03169_));
 sky130_fd_sc_hd__a22oi_4 _17875_ (.A1(\CPU_Xreg_value_a4[16][11] ),
    .A2(_02979_),
    .B1(\CPU_Xreg_value_a4[30][11] ),
    .B2(_02980_),
    .Y(_03170_));
 sky130_fd_sc_hd__o22a_4 _17876_ (.A1(_02017_),
    .A2(_02982_),
    .B1(_02002_),
    .B2(_02983_),
    .X(_03171_));
 sky130_fd_sc_hd__o22a_4 _17877_ (.A1(_02015_),
    .A2(_02985_),
    .B1(_02018_),
    .B2(_02986_),
    .X(_03172_));
 sky130_fd_sc_hd__and4_4 _17878_ (.A(_03169_),
    .B(_03170_),
    .C(_03171_),
    .D(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__inv_2 _17879_ (.A(\CPU_Xreg_value_a4[26][11] ),
    .Y(_03174_));
 sky130_fd_sc_hd__o22a_4 _17880_ (.A1(_03174_),
    .A2(_02990_),
    .B1(_02003_),
    .B2(_02991_),
    .X(_03175_));
 sky130_fd_sc_hd__o22a_4 _17881_ (.A1(_02020_),
    .A2(_02993_),
    .B1(_02009_),
    .B2(_02994_),
    .X(_03176_));
 sky130_fd_sc_hd__a22oi_4 _17882_ (.A1(\CPU_Xreg_value_a4[23][11] ),
    .A2(_02996_),
    .B1(\CPU_Xreg_value_a4[31][11] ),
    .B2(_02997_),
    .Y(_03177_));
 sky130_fd_sc_hd__inv_2 _17883_ (.A(\CPU_Xreg_value_a4[19][11] ),
    .Y(_03178_));
 sky130_fd_sc_hd__o22a_4 _17884_ (.A1(_03178_),
    .A2(_03000_),
    .B1(_02024_),
    .B2(_03001_),
    .X(_03179_));
 sky130_fd_sc_hd__and4_4 _17885_ (.A(_03175_),
    .B(_03176_),
    .C(_03177_),
    .D(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__o22a_4 _17886_ (.A1(_02000_),
    .A2(_03004_),
    .B1(_02023_),
    .B2(_03005_),
    .X(_03181_));
 sky130_fd_sc_hd__inv_2 _17887_ (.A(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__inv_2 _17888_ (.A(\CPU_Xreg_value_a4[25][11] ),
    .Y(_03183_));
 sky130_fd_sc_hd__a2bb2o_4 _17889_ (.A1_N(_03183_),
    .A2_N(_03009_),
    .B1(\CPU_Xreg_value_a4[24][11] ),
    .B2(_03010_),
    .X(_03184_));
 sky130_fd_sc_hd__inv_2 _17890_ (.A(\CPU_Xreg_value_a4[17][11] ),
    .Y(_03185_));
 sky130_fd_sc_hd__a2bb2o_4 _17891_ (.A1_N(_03185_),
    .A2_N(_03014_),
    .B1(\CPU_Xreg_value_a4[22][11] ),
    .B2(_03015_),
    .X(_03186_));
 sky130_fd_sc_hd__a211o_4 _17892_ (.A1(\CPU_Xreg_value_a4[13][11] ),
    .A2(_03012_),
    .B1(_03152_),
    .C1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__inv_2 _17893_ (.A(\CPU_Xreg_value_a4[18][11] ),
    .Y(_03188_));
 sky130_fd_sc_hd__a2bb2o_4 _17894_ (.A1_N(_03188_),
    .A2_N(_03019_),
    .B1(\CPU_Xreg_value_a4[28][11] ),
    .B2(_03020_),
    .X(_03189_));
 sky130_fd_sc_hd__o22a_4 _17895_ (.A1(_02006_),
    .A2(_03022_),
    .B1(_02014_),
    .B2(_03023_),
    .X(_03190_));
 sky130_fd_sc_hd__inv_2 _17896_ (.A(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__inv_2 _17897_ (.A(\CPU_Xreg_value_a4[21][11] ),
    .Y(_03192_));
 sky130_fd_sc_hd__a2bb2o_4 _17898_ (.A1_N(_03192_),
    .A2_N(_03027_),
    .B1(\CPU_Xreg_value_a4[20][11] ),
    .B2(_03028_),
    .X(_03193_));
 sky130_fd_sc_hd__inv_2 _17899_ (.A(\CPU_Xreg_value_a4[27][11] ),
    .Y(_03194_));
 sky130_fd_sc_hd__a2bb2o_4 _17900_ (.A1_N(_03194_),
    .A2_N(_03031_),
    .B1(\CPU_Xreg_value_a4[29][11] ),
    .B2(_03032_),
    .X(_03195_));
 sky130_fd_sc_hd__or4_4 _17901_ (.A(_03189_),
    .B(_03191_),
    .C(_03193_),
    .D(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__or4_4 _17902_ (.A(_03182_),
    .B(_03184_),
    .C(_03187_),
    .D(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__inv_2 _17903_ (.A(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__a32o_4 _17904_ (.A1(_03173_),
    .A2(_03180_),
    .A3(_03198_),
    .B1(_06129_),
    .B2(_03037_),
    .X(_03199_));
 sky130_fd_sc_hd__inv_2 _17905_ (.A(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o22a_4 _17906_ (.A1(_06768_),
    .A2(_02974_),
    .B1(_02975_),
    .B2(_03200_),
    .X(\CPU_src2_value_a2[11] ));
 sky130_fd_sc_hd__buf_2 _17907_ (.A(_02669_),
    .X(_03201_));
 sky130_fd_sc_hd__buf_2 _17908_ (.A(_02672_),
    .X(_03202_));
 sky130_fd_sc_hd__buf_2 _17909_ (.A(_02681_),
    .X(_03203_));
 sky130_fd_sc_hd__buf_2 _17910_ (.A(_02686_),
    .X(_03204_));
 sky130_fd_sc_hd__o22a_4 _17911_ (.A1(_02043_),
    .A2(_03203_),
    .B1(_02060_),
    .B2(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__buf_2 _17912_ (.A(_02693_),
    .X(_03206_));
 sky130_fd_sc_hd__buf_2 _17913_ (.A(_02699_),
    .X(_03207_));
 sky130_fd_sc_hd__a22oi_4 _17914_ (.A1(\CPU_Xreg_value_a4[16][12] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][12] ),
    .B2(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__buf_2 _17915_ (.A(_02704_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_2 _17916_ (.A(_02708_),
    .X(_03210_));
 sky130_fd_sc_hd__o22a_4 _17917_ (.A1(_02053_),
    .A2(_03209_),
    .B1(_02033_),
    .B2(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__buf_2 _17918_ (.A(_02712_),
    .X(_03212_));
 sky130_fd_sc_hd__buf_2 _17919_ (.A(_02715_),
    .X(_03213_));
 sky130_fd_sc_hd__o22a_4 _17920_ (.A1(_02050_),
    .A2(_03212_),
    .B1(_02055_),
    .B2(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__and4_4 _17921_ (.A(_03205_),
    .B(_03208_),
    .C(_03211_),
    .D(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__inv_2 _17922_ (.A(\CPU_Xreg_value_a4[26][12] ),
    .Y(_03216_));
 sky130_fd_sc_hd__buf_2 _17923_ (.A(_02721_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_2 _17924_ (.A(_02724_),
    .X(_03218_));
 sky130_fd_sc_hd__o22a_4 _17925_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_02035_),
    .B2(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__buf_2 _17926_ (.A(_02728_),
    .X(_03220_));
 sky130_fd_sc_hd__buf_2 _17927_ (.A(_02731_),
    .X(_03221_));
 sky130_fd_sc_hd__o22a_4 _17928_ (.A1(_02058_),
    .A2(_03220_),
    .B1(_02041_),
    .B2(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__buf_2 _17929_ (.A(_02736_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_2 _17930_ (.A(_02740_),
    .X(_03224_));
 sky130_fd_sc_hd__a22oi_4 _17931_ (.A1(\CPU_Xreg_value_a4[23][12] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][12] ),
    .B2(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__inv_2 _17932_ (.A(\CPU_Xreg_value_a4[19][12] ),
    .Y(_03226_));
 sky130_fd_sc_hd__buf_2 _17933_ (.A(_02744_),
    .X(_03227_));
 sky130_fd_sc_hd__buf_2 _17934_ (.A(_02747_),
    .X(_03228_));
 sky130_fd_sc_hd__o22a_4 _17935_ (.A1(_03226_),
    .A2(_03227_),
    .B1(_02065_),
    .B2(_03228_),
    .X(_03229_));
 sky130_fd_sc_hd__and4_4 _17936_ (.A(_03219_),
    .B(_03222_),
    .C(_03225_),
    .D(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__buf_2 _17937_ (.A(_02752_),
    .X(_03231_));
 sky130_fd_sc_hd__buf_2 _17938_ (.A(_02756_),
    .X(_03232_));
 sky130_fd_sc_hd__o22a_4 _17939_ (.A1(_02031_),
    .A2(_03231_),
    .B1(_02063_),
    .B2(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__inv_2 _17940_ (.A(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__inv_2 _17941_ (.A(\CPU_Xreg_value_a4[25][12] ),
    .Y(_03235_));
 sky130_fd_sc_hd__buf_2 _17942_ (.A(_02761_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_2 _17943_ (.A(_02765_),
    .X(_03237_));
 sky130_fd_sc_hd__a2bb2o_4 _17944_ (.A1_N(_03235_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][12] ),
    .B2(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_2 _17945_ (.A(_02771_),
    .X(_03239_));
 sky130_fd_sc_hd__inv_2 _17946_ (.A(\CPU_Xreg_value_a4[17][12] ),
    .Y(_03240_));
 sky130_fd_sc_hd__buf_2 _17947_ (.A(_02778_),
    .X(_03241_));
 sky130_fd_sc_hd__buf_2 _17948_ (.A(_02783_),
    .X(_03242_));
 sky130_fd_sc_hd__a2bb2o_4 _17949_ (.A1_N(_03240_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][12] ),
    .B2(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__a211o_4 _17950_ (.A1(\CPU_Xreg_value_a4[13][12] ),
    .A2(_03239_),
    .B1(_03152_),
    .C1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__inv_2 _17951_ (.A(\CPU_Xreg_value_a4[18][12] ),
    .Y(_03245_));
 sky130_fd_sc_hd__buf_2 _17952_ (.A(_02789_),
    .X(_03246_));
 sky130_fd_sc_hd__buf_2 _17953_ (.A(_02793_),
    .X(_03247_));
 sky130_fd_sc_hd__a2bb2o_4 _17954_ (.A1_N(_03245_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][12] ),
    .B2(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_2 _17955_ (.A(_02797_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_2 _17956_ (.A(_02800_),
    .X(_03250_));
 sky130_fd_sc_hd__o22a_4 _17957_ (.A1(_02039_),
    .A2(_03249_),
    .B1(_02048_),
    .B2(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__inv_2 _17958_ (.A(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__inv_2 _17959_ (.A(\CPU_Xreg_value_a4[21][12] ),
    .Y(_03253_));
 sky130_fd_sc_hd__buf_2 _17960_ (.A(_02805_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_2 _17961_ (.A(_02809_),
    .X(_03255_));
 sky130_fd_sc_hd__a2bb2o_4 _17962_ (.A1_N(_03253_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][12] ),
    .B2(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__inv_2 _17963_ (.A(\CPU_Xreg_value_a4[27][12] ),
    .Y(_03257_));
 sky130_fd_sc_hd__buf_2 _17964_ (.A(_02813_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_2 _17965_ (.A(_02817_),
    .X(_03259_));
 sky130_fd_sc_hd__a2bb2o_4 _17966_ (.A1_N(_03257_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][12] ),
    .B2(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__or4_4 _17967_ (.A(_03248_),
    .B(_03252_),
    .C(_03256_),
    .D(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__or4_4 _17968_ (.A(_03234_),
    .B(_03238_),
    .C(_03244_),
    .D(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__inv_2 _17969_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__buf_2 _17970_ (.A(_02823_),
    .X(_03264_));
 sky130_fd_sc_hd__a32o_4 _17971_ (.A1(_03215_),
    .A2(_03230_),
    .A3(_03263_),
    .B1(_06128_),
    .B2(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__inv_2 _17972_ (.A(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o22a_4 _17973_ (.A1(_06750_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03266_),
    .X(\CPU_src2_value_a2[12] ));
 sky130_fd_sc_hd__o22a_4 _17974_ (.A1(_02084_),
    .A2(_03203_),
    .B1(_02095_),
    .B2(_03204_),
    .X(_03267_));
 sky130_fd_sc_hd__a22oi_4 _17975_ (.A1(\CPU_Xreg_value_a4[16][13] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][13] ),
    .B2(_03207_),
    .Y(_03268_));
 sky130_fd_sc_hd__o22a_4 _17976_ (.A1(_02091_),
    .A2(_03209_),
    .B1(_02076_),
    .B2(_03210_),
    .X(_03269_));
 sky130_fd_sc_hd__o22a_4 _17977_ (.A1(_02089_),
    .A2(_03212_),
    .B1(_02092_),
    .B2(_03213_),
    .X(_03270_));
 sky130_fd_sc_hd__and4_4 _17978_ (.A(_03267_),
    .B(_03268_),
    .C(_03269_),
    .D(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__inv_2 _17979_ (.A(\CPU_Xreg_value_a4[26][13] ),
    .Y(_03272_));
 sky130_fd_sc_hd__o22a_4 _17980_ (.A1(_03272_),
    .A2(_03217_),
    .B1(_02077_),
    .B2(_03218_),
    .X(_03273_));
 sky130_fd_sc_hd__o22a_4 _17981_ (.A1(_02094_),
    .A2(_03220_),
    .B1(_02083_),
    .B2(_03221_),
    .X(_03274_));
 sky130_fd_sc_hd__a22oi_4 _17982_ (.A1(\CPU_Xreg_value_a4[23][13] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][13] ),
    .B2(_03224_),
    .Y(_03275_));
 sky130_fd_sc_hd__inv_2 _17983_ (.A(\CPU_Xreg_value_a4[19][13] ),
    .Y(_03276_));
 sky130_fd_sc_hd__o22a_4 _17984_ (.A1(_03276_),
    .A2(_03227_),
    .B1(_02098_),
    .B2(_03228_),
    .X(_03277_));
 sky130_fd_sc_hd__and4_4 _17985_ (.A(_03273_),
    .B(_03274_),
    .C(_03275_),
    .D(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__o22a_4 _17986_ (.A1(_02072_),
    .A2(_03231_),
    .B1(_02097_),
    .B2(_03232_),
    .X(_03279_));
 sky130_fd_sc_hd__inv_2 _17987_ (.A(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__inv_2 _17988_ (.A(\CPU_Xreg_value_a4[25][13] ),
    .Y(_03281_));
 sky130_fd_sc_hd__a2bb2o_4 _17989_ (.A1_N(_03281_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][13] ),
    .B2(_03237_),
    .X(_03282_));
 sky130_fd_sc_hd__inv_2 _17990_ (.A(\CPU_Xreg_value_a4[17][13] ),
    .Y(_03283_));
 sky130_fd_sc_hd__a2bb2o_4 _17991_ (.A1_N(_03283_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][13] ),
    .B2(_03242_),
    .X(_03284_));
 sky130_fd_sc_hd__a211o_4 _17992_ (.A1(\CPU_Xreg_value_a4[13][13] ),
    .A2(_03239_),
    .B1(_03152_),
    .C1(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__inv_2 _17993_ (.A(\CPU_Xreg_value_a4[18][13] ),
    .Y(_03286_));
 sky130_fd_sc_hd__a2bb2o_4 _17994_ (.A1_N(_03286_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][13] ),
    .B2(_03247_),
    .X(_03287_));
 sky130_fd_sc_hd__o22a_4 _17995_ (.A1(_02080_),
    .A2(_03249_),
    .B1(_02088_),
    .B2(_03250_),
    .X(_03288_));
 sky130_fd_sc_hd__inv_2 _17996_ (.A(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__inv_2 _17997_ (.A(\CPU_Xreg_value_a4[21][13] ),
    .Y(_03290_));
 sky130_fd_sc_hd__a2bb2o_4 _17998_ (.A1_N(_03290_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][13] ),
    .B2(_03255_),
    .X(_03291_));
 sky130_fd_sc_hd__inv_2 _17999_ (.A(\CPU_Xreg_value_a4[27][13] ),
    .Y(_03292_));
 sky130_fd_sc_hd__a2bb2o_4 _18000_ (.A1_N(_03292_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][13] ),
    .B2(_03259_),
    .X(_03293_));
 sky130_fd_sc_hd__or4_4 _18001_ (.A(_03287_),
    .B(_03289_),
    .C(_03291_),
    .D(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__or4_4 _18002_ (.A(_03280_),
    .B(_03282_),
    .C(_03285_),
    .D(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__inv_2 _18003_ (.A(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__a32o_4 _18004_ (.A1(_03271_),
    .A2(_03278_),
    .A3(_03296_),
    .B1(_06127_),
    .B2(_03264_),
    .X(_03297_));
 sky130_fd_sc_hd__inv_2 _18005_ (.A(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__o22a_4 _18006_ (.A1(_06741_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03298_),
    .X(\CPU_src2_value_a2[13] ));
 sky130_fd_sc_hd__o22a_4 _18007_ (.A1(_02112_),
    .A2(_03203_),
    .B1(_02123_),
    .B2(_03204_),
    .X(_03299_));
 sky130_fd_sc_hd__a22oi_4 _18008_ (.A1(\CPU_Xreg_value_a4[16][14] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][14] ),
    .B2(_03207_),
    .Y(_03300_));
 sky130_fd_sc_hd__o22a_4 _18009_ (.A1(_02119_),
    .A2(_03209_),
    .B1(_02105_),
    .B2(_03210_),
    .X(_03301_));
 sky130_fd_sc_hd__o22a_4 _18010_ (.A1(_02117_),
    .A2(_03212_),
    .B1(_02120_),
    .B2(_03213_),
    .X(_03302_));
 sky130_fd_sc_hd__and4_4 _18011_ (.A(_03299_),
    .B(_03300_),
    .C(_03301_),
    .D(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__inv_2 _18012_ (.A(\CPU_Xreg_value_a4[26][14] ),
    .Y(_03304_));
 sky130_fd_sc_hd__o22a_4 _18013_ (.A1(_03304_),
    .A2(_03217_),
    .B1(_02106_),
    .B2(_03218_),
    .X(_03305_));
 sky130_fd_sc_hd__o22a_4 _18014_ (.A1(_02122_),
    .A2(_03220_),
    .B1(_02111_),
    .B2(_03221_),
    .X(_03306_));
 sky130_fd_sc_hd__a22oi_4 _18015_ (.A1(\CPU_Xreg_value_a4[23][14] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][14] ),
    .B2(_03224_),
    .Y(_03307_));
 sky130_fd_sc_hd__inv_2 _18016_ (.A(\CPU_Xreg_value_a4[19][14] ),
    .Y(_03308_));
 sky130_fd_sc_hd__o22a_4 _18017_ (.A1(_03308_),
    .A2(_03227_),
    .B1(_02126_),
    .B2(_03228_),
    .X(_03309_));
 sky130_fd_sc_hd__and4_4 _18018_ (.A(_03305_),
    .B(_03306_),
    .C(_03307_),
    .D(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__o22a_4 _18019_ (.A1(_02103_),
    .A2(_03231_),
    .B1(_02125_),
    .B2(_03232_),
    .X(_03311_));
 sky130_fd_sc_hd__inv_2 _18020_ (.A(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__inv_2 _18021_ (.A(\CPU_Xreg_value_a4[25][14] ),
    .Y(_03313_));
 sky130_fd_sc_hd__a2bb2o_4 _18022_ (.A1_N(_03313_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][14] ),
    .B2(_03237_),
    .X(_03314_));
 sky130_fd_sc_hd__inv_2 _18023_ (.A(\CPU_Xreg_value_a4[17][14] ),
    .Y(_03315_));
 sky130_fd_sc_hd__a2bb2o_4 _18024_ (.A1_N(_03315_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][14] ),
    .B2(_03242_),
    .X(_03316_));
 sky130_fd_sc_hd__a211o_4 _18025_ (.A1(\CPU_Xreg_value_a4[13][14] ),
    .A2(_03239_),
    .B1(_03152_),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__inv_2 _18026_ (.A(\CPU_Xreg_value_a4[18][14] ),
    .Y(_03318_));
 sky130_fd_sc_hd__a2bb2o_4 _18027_ (.A1_N(_03318_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][14] ),
    .B2(_03247_),
    .X(_03319_));
 sky130_fd_sc_hd__o22a_4 _18028_ (.A1(_02109_),
    .A2(_03249_),
    .B1(_02116_),
    .B2(_03250_),
    .X(_03320_));
 sky130_fd_sc_hd__inv_2 _18029_ (.A(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__inv_2 _18030_ (.A(\CPU_Xreg_value_a4[21][14] ),
    .Y(_03322_));
 sky130_fd_sc_hd__a2bb2o_4 _18031_ (.A1_N(_03322_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][14] ),
    .B2(_03255_),
    .X(_03323_));
 sky130_fd_sc_hd__inv_2 _18032_ (.A(\CPU_Xreg_value_a4[27][14] ),
    .Y(_03324_));
 sky130_fd_sc_hd__a2bb2o_4 _18033_ (.A1_N(_03324_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][14] ),
    .B2(_03259_),
    .X(_03325_));
 sky130_fd_sc_hd__or4_4 _18034_ (.A(_03319_),
    .B(_03321_),
    .C(_03323_),
    .D(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__or4_4 _18035_ (.A(_03312_),
    .B(_03314_),
    .C(_03317_),
    .D(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__inv_2 _18036_ (.A(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__a32o_4 _18037_ (.A1(_03303_),
    .A2(_03310_),
    .A3(_03328_),
    .B1(_06125_),
    .B2(_03264_),
    .X(_03329_));
 sky130_fd_sc_hd__inv_2 _18038_ (.A(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__o22a_4 _18039_ (.A1(_06731_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03330_),
    .X(\CPU_src2_value_a2[14] ));
 sky130_fd_sc_hd__o22a_4 _18040_ (.A1(_02140_),
    .A2(_03203_),
    .B1(_02151_),
    .B2(_03204_),
    .X(_03331_));
 sky130_fd_sc_hd__a22oi_4 _18041_ (.A1(\CPU_Xreg_value_a4[16][15] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][15] ),
    .B2(_03207_),
    .Y(_03332_));
 sky130_fd_sc_hd__o22a_4 _18042_ (.A1(_02147_),
    .A2(_03209_),
    .B1(_02133_),
    .B2(_03210_),
    .X(_03333_));
 sky130_fd_sc_hd__o22a_4 _18043_ (.A1(_02145_),
    .A2(_03212_),
    .B1(_02148_),
    .B2(_03213_),
    .X(_03334_));
 sky130_fd_sc_hd__and4_4 _18044_ (.A(_03331_),
    .B(_03332_),
    .C(_03333_),
    .D(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__inv_2 _18045_ (.A(\CPU_Xreg_value_a4[26][15] ),
    .Y(_03336_));
 sky130_fd_sc_hd__o22a_4 _18046_ (.A1(_03336_),
    .A2(_03217_),
    .B1(_02134_),
    .B2(_03218_),
    .X(_03337_));
 sky130_fd_sc_hd__o22a_4 _18047_ (.A1(_02150_),
    .A2(_03220_),
    .B1(_02139_),
    .B2(_03221_),
    .X(_03338_));
 sky130_fd_sc_hd__a22oi_4 _18048_ (.A1(\CPU_Xreg_value_a4[23][15] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][15] ),
    .B2(_03224_),
    .Y(_03339_));
 sky130_fd_sc_hd__inv_2 _18049_ (.A(\CPU_Xreg_value_a4[19][15] ),
    .Y(_03340_));
 sky130_fd_sc_hd__o22a_4 _18050_ (.A1(_03340_),
    .A2(_03227_),
    .B1(_02154_),
    .B2(_03228_),
    .X(_03341_));
 sky130_fd_sc_hd__and4_4 _18051_ (.A(_03337_),
    .B(_03338_),
    .C(_03339_),
    .D(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__o22a_4 _18052_ (.A1(_02131_),
    .A2(_03231_),
    .B1(_02153_),
    .B2(_03232_),
    .X(_03343_));
 sky130_fd_sc_hd__inv_2 _18053_ (.A(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__inv_2 _18054_ (.A(\CPU_Xreg_value_a4[25][15] ),
    .Y(_03345_));
 sky130_fd_sc_hd__a2bb2o_4 _18055_ (.A1_N(_03345_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][15] ),
    .B2(_03237_),
    .X(_03346_));
 sky130_fd_sc_hd__inv_2 _18056_ (.A(\CPU_Xreg_value_a4[17][15] ),
    .Y(_03347_));
 sky130_fd_sc_hd__a2bb2o_4 _18057_ (.A1_N(_03347_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][15] ),
    .B2(_03242_),
    .X(_03348_));
 sky130_fd_sc_hd__a211o_4 _18058_ (.A1(\CPU_Xreg_value_a4[13][15] ),
    .A2(_03239_),
    .B1(_03152_),
    .C1(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__inv_2 _18059_ (.A(\CPU_Xreg_value_a4[18][15] ),
    .Y(_03350_));
 sky130_fd_sc_hd__a2bb2o_4 _18060_ (.A1_N(_03350_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][15] ),
    .B2(_03247_),
    .X(_03351_));
 sky130_fd_sc_hd__o22a_4 _18061_ (.A1(_02137_),
    .A2(_03249_),
    .B1(_02144_),
    .B2(_03250_),
    .X(_03352_));
 sky130_fd_sc_hd__inv_2 _18062_ (.A(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__inv_2 _18063_ (.A(\CPU_Xreg_value_a4[21][15] ),
    .Y(_03354_));
 sky130_fd_sc_hd__a2bb2o_4 _18064_ (.A1_N(_03354_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][15] ),
    .B2(_03255_),
    .X(_03355_));
 sky130_fd_sc_hd__inv_2 _18065_ (.A(\CPU_Xreg_value_a4[27][15] ),
    .Y(_03356_));
 sky130_fd_sc_hd__a2bb2o_4 _18066_ (.A1_N(_03356_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][15] ),
    .B2(_03259_),
    .X(_03357_));
 sky130_fd_sc_hd__or4_4 _18067_ (.A(_03351_),
    .B(_03353_),
    .C(_03355_),
    .D(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__or4_4 _18068_ (.A(_03344_),
    .B(_03346_),
    .C(_03349_),
    .D(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__inv_2 _18069_ (.A(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__a32o_4 _18070_ (.A1(_03335_),
    .A2(_03342_),
    .A3(_03360_),
    .B1(_06124_),
    .B2(_03264_),
    .X(_03361_));
 sky130_fd_sc_hd__inv_2 _18071_ (.A(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__o22a_4 _18072_ (.A1(_06722_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03362_),
    .X(\CPU_src2_value_a2[15] ));
 sky130_fd_sc_hd__o22a_4 _18073_ (.A1(_02168_),
    .A2(_03203_),
    .B1(_02179_),
    .B2(_03204_),
    .X(_03363_));
 sky130_fd_sc_hd__a22oi_4 _18074_ (.A1(\CPU_Xreg_value_a4[16][16] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][16] ),
    .B2(_03207_),
    .Y(_03364_));
 sky130_fd_sc_hd__o22a_4 _18075_ (.A1(_02175_),
    .A2(_03209_),
    .B1(_02161_),
    .B2(_03210_),
    .X(_03365_));
 sky130_fd_sc_hd__o22a_4 _18076_ (.A1(_02173_),
    .A2(_03212_),
    .B1(_02176_),
    .B2(_03213_),
    .X(_03366_));
 sky130_fd_sc_hd__and4_4 _18077_ (.A(_03363_),
    .B(_03364_),
    .C(_03365_),
    .D(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__inv_2 _18078_ (.A(\CPU_Xreg_value_a4[26][16] ),
    .Y(_03368_));
 sky130_fd_sc_hd__o22a_4 _18079_ (.A1(_03368_),
    .A2(_03217_),
    .B1(_02162_),
    .B2(_03218_),
    .X(_03369_));
 sky130_fd_sc_hd__o22a_4 _18080_ (.A1(_02178_),
    .A2(_03220_),
    .B1(_02167_),
    .B2(_03221_),
    .X(_03370_));
 sky130_fd_sc_hd__a22oi_4 _18081_ (.A1(\CPU_Xreg_value_a4[23][16] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][16] ),
    .B2(_03224_),
    .Y(_03371_));
 sky130_fd_sc_hd__inv_2 _18082_ (.A(\CPU_Xreg_value_a4[19][16] ),
    .Y(_03372_));
 sky130_fd_sc_hd__o22a_4 _18083_ (.A1(_03372_),
    .A2(_03227_),
    .B1(_02182_),
    .B2(_03228_),
    .X(_03373_));
 sky130_fd_sc_hd__and4_4 _18084_ (.A(_03369_),
    .B(_03370_),
    .C(_03371_),
    .D(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__o22a_4 _18085_ (.A1(_02159_),
    .A2(_03231_),
    .B1(_02181_),
    .B2(_03232_),
    .X(_03375_));
 sky130_fd_sc_hd__inv_2 _18086_ (.A(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__inv_2 _18087_ (.A(\CPU_Xreg_value_a4[25][16] ),
    .Y(_03377_));
 sky130_fd_sc_hd__a2bb2o_4 _18088_ (.A1_N(_03377_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][16] ),
    .B2(_03237_),
    .X(_03378_));
 sky130_fd_sc_hd__buf_2 _18089_ (.A(_02774_),
    .X(_03379_));
 sky130_fd_sc_hd__inv_2 _18090_ (.A(\CPU_Xreg_value_a4[17][16] ),
    .Y(_03380_));
 sky130_fd_sc_hd__a2bb2o_4 _18091_ (.A1_N(_03380_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][16] ),
    .B2(_03242_),
    .X(_03381_));
 sky130_fd_sc_hd__a211o_4 _18092_ (.A1(\CPU_Xreg_value_a4[13][16] ),
    .A2(_03239_),
    .B1(_03379_),
    .C1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__inv_2 _18093_ (.A(\CPU_Xreg_value_a4[18][16] ),
    .Y(_03383_));
 sky130_fd_sc_hd__a2bb2o_4 _18094_ (.A1_N(_03383_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][16] ),
    .B2(_03247_),
    .X(_03384_));
 sky130_fd_sc_hd__o22a_4 _18095_ (.A1(_02165_),
    .A2(_03249_),
    .B1(_02172_),
    .B2(_03250_),
    .X(_03385_));
 sky130_fd_sc_hd__inv_2 _18096_ (.A(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__inv_2 _18097_ (.A(\CPU_Xreg_value_a4[21][16] ),
    .Y(_03387_));
 sky130_fd_sc_hd__a2bb2o_4 _18098_ (.A1_N(_03387_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][16] ),
    .B2(_03255_),
    .X(_03388_));
 sky130_fd_sc_hd__inv_2 _18099_ (.A(\CPU_Xreg_value_a4[27][16] ),
    .Y(_03389_));
 sky130_fd_sc_hd__a2bb2o_4 _18100_ (.A1_N(_03389_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][16] ),
    .B2(_03259_),
    .X(_03390_));
 sky130_fd_sc_hd__or4_4 _18101_ (.A(_03384_),
    .B(_03386_),
    .C(_03388_),
    .D(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__or4_4 _18102_ (.A(_03376_),
    .B(_03378_),
    .C(_03382_),
    .D(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__inv_2 _18103_ (.A(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__a32o_4 _18104_ (.A1(_03367_),
    .A2(_03374_),
    .A3(_03393_),
    .B1(_06123_),
    .B2(_03264_),
    .X(_03394_));
 sky130_fd_sc_hd__inv_2 _18105_ (.A(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__o22a_4 _18106_ (.A1(_06699_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03395_),
    .X(\CPU_src2_value_a2[16] ));
 sky130_fd_sc_hd__o22a_4 _18107_ (.A1(_02197_),
    .A2(_03203_),
    .B1(_02208_),
    .B2(_03204_),
    .X(_03396_));
 sky130_fd_sc_hd__a22oi_4 _18108_ (.A1(\CPU_Xreg_value_a4[16][17] ),
    .A2(_03206_),
    .B1(\CPU_Xreg_value_a4[30][17] ),
    .B2(_03207_),
    .Y(_03397_));
 sky130_fd_sc_hd__o22a_4 _18109_ (.A1(_02204_),
    .A2(_03209_),
    .B1(_02189_),
    .B2(_03210_),
    .X(_03398_));
 sky130_fd_sc_hd__o22a_4 _18110_ (.A1(_02202_),
    .A2(_03212_),
    .B1(_02205_),
    .B2(_03213_),
    .X(_03399_));
 sky130_fd_sc_hd__and4_4 _18111_ (.A(_03396_),
    .B(_03397_),
    .C(_03398_),
    .D(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__inv_2 _18112_ (.A(\CPU_Xreg_value_a4[26][17] ),
    .Y(_03401_));
 sky130_fd_sc_hd__o22a_4 _18113_ (.A1(_03401_),
    .A2(_03217_),
    .B1(_02190_),
    .B2(_03218_),
    .X(_03402_));
 sky130_fd_sc_hd__o22a_4 _18114_ (.A1(_02207_),
    .A2(_03220_),
    .B1(_02196_),
    .B2(_03221_),
    .X(_03403_));
 sky130_fd_sc_hd__a22oi_4 _18115_ (.A1(\CPU_Xreg_value_a4[23][17] ),
    .A2(_03223_),
    .B1(\CPU_Xreg_value_a4[31][17] ),
    .B2(_03224_),
    .Y(_03404_));
 sky130_fd_sc_hd__inv_2 _18116_ (.A(\CPU_Xreg_value_a4[19][17] ),
    .Y(_03405_));
 sky130_fd_sc_hd__o22a_4 _18117_ (.A1(_03405_),
    .A2(_03227_),
    .B1(_02211_),
    .B2(_03228_),
    .X(_03406_));
 sky130_fd_sc_hd__and4_4 _18118_ (.A(_03402_),
    .B(_03403_),
    .C(_03404_),
    .D(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__o22a_4 _18119_ (.A1(_02187_),
    .A2(_03231_),
    .B1(_02210_),
    .B2(_03232_),
    .X(_03408_));
 sky130_fd_sc_hd__inv_2 _18120_ (.A(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__inv_2 _18121_ (.A(\CPU_Xreg_value_a4[25][17] ),
    .Y(_03410_));
 sky130_fd_sc_hd__a2bb2o_4 _18122_ (.A1_N(_03410_),
    .A2_N(_03236_),
    .B1(\CPU_Xreg_value_a4[24][17] ),
    .B2(_03237_),
    .X(_03411_));
 sky130_fd_sc_hd__inv_2 _18123_ (.A(\CPU_Xreg_value_a4[17][17] ),
    .Y(_03412_));
 sky130_fd_sc_hd__a2bb2o_4 _18124_ (.A1_N(_03412_),
    .A2_N(_03241_),
    .B1(\CPU_Xreg_value_a4[22][17] ),
    .B2(_03242_),
    .X(_03413_));
 sky130_fd_sc_hd__a211o_4 _18125_ (.A1(\CPU_Xreg_value_a4[13][17] ),
    .A2(_03239_),
    .B1(_03379_),
    .C1(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__inv_2 _18126_ (.A(\CPU_Xreg_value_a4[18][17] ),
    .Y(_03415_));
 sky130_fd_sc_hd__a2bb2o_4 _18127_ (.A1_N(_03415_),
    .A2_N(_03246_),
    .B1(\CPU_Xreg_value_a4[28][17] ),
    .B2(_03247_),
    .X(_03416_));
 sky130_fd_sc_hd__o22a_4 _18128_ (.A1(_02193_),
    .A2(_03249_),
    .B1(_02201_),
    .B2(_03250_),
    .X(_03417_));
 sky130_fd_sc_hd__inv_2 _18129_ (.A(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__inv_2 _18130_ (.A(\CPU_Xreg_value_a4[21][17] ),
    .Y(_03419_));
 sky130_fd_sc_hd__a2bb2o_4 _18131_ (.A1_N(_03419_),
    .A2_N(_03254_),
    .B1(\CPU_Xreg_value_a4[20][17] ),
    .B2(_03255_),
    .X(_03420_));
 sky130_fd_sc_hd__inv_2 _18132_ (.A(\CPU_Xreg_value_a4[27][17] ),
    .Y(_03421_));
 sky130_fd_sc_hd__a2bb2o_4 _18133_ (.A1_N(_03421_),
    .A2_N(_03258_),
    .B1(\CPU_Xreg_value_a4[29][17] ),
    .B2(_03259_),
    .X(_03422_));
 sky130_fd_sc_hd__or4_4 _18134_ (.A(_03416_),
    .B(_03418_),
    .C(_03420_),
    .D(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__or4_4 _18135_ (.A(_03409_),
    .B(_03411_),
    .C(_03414_),
    .D(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__inv_2 _18136_ (.A(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__a32o_4 _18137_ (.A1(_03400_),
    .A2(_03407_),
    .A3(_03425_),
    .B1(_06122_),
    .B2(_03264_),
    .X(_03426_));
 sky130_fd_sc_hd__inv_2 _18138_ (.A(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__o22a_4 _18139_ (.A1(_06690_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03427_),
    .X(\CPU_src2_value_a2[17] ));
 sky130_fd_sc_hd__buf_2 _18140_ (.A(_02669_),
    .X(_03428_));
 sky130_fd_sc_hd__buf_2 _18141_ (.A(_02672_),
    .X(_03429_));
 sky130_fd_sc_hd__buf_2 _18142_ (.A(_02681_),
    .X(_03430_));
 sky130_fd_sc_hd__buf_2 _18143_ (.A(_02686_),
    .X(_03431_));
 sky130_fd_sc_hd__o22a_4 _18144_ (.A1(_02230_),
    .A2(_03430_),
    .B1(_02247_),
    .B2(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__buf_2 _18145_ (.A(_02693_),
    .X(_03433_));
 sky130_fd_sc_hd__buf_2 _18146_ (.A(_02699_),
    .X(_03434_));
 sky130_fd_sc_hd__a22oi_4 _18147_ (.A1(\CPU_Xreg_value_a4[16][18] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][18] ),
    .B2(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__buf_2 _18148_ (.A(_02704_),
    .X(_03436_));
 sky130_fd_sc_hd__buf_2 _18149_ (.A(_02708_),
    .X(_03437_));
 sky130_fd_sc_hd__o22a_4 _18150_ (.A1(_02240_),
    .A2(_03436_),
    .B1(_02220_),
    .B2(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__buf_2 _18151_ (.A(_02712_),
    .X(_03439_));
 sky130_fd_sc_hd__buf_2 _18152_ (.A(_02715_),
    .X(_03440_));
 sky130_fd_sc_hd__o22a_4 _18153_ (.A1(_02237_),
    .A2(_03439_),
    .B1(_02242_),
    .B2(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__and4_4 _18154_ (.A(_03432_),
    .B(_03435_),
    .C(_03438_),
    .D(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__inv_2 _18155_ (.A(\CPU_Xreg_value_a4[26][18] ),
    .Y(_03443_));
 sky130_fd_sc_hd__buf_2 _18156_ (.A(_02721_),
    .X(_03444_));
 sky130_fd_sc_hd__buf_2 _18157_ (.A(_02724_),
    .X(_03445_));
 sky130_fd_sc_hd__o22a_4 _18158_ (.A1(_03443_),
    .A2(_03444_),
    .B1(_02222_),
    .B2(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__buf_2 _18159_ (.A(_02728_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_2 _18160_ (.A(_02731_),
    .X(_03448_));
 sky130_fd_sc_hd__o22a_4 _18161_ (.A1(_02245_),
    .A2(_03447_),
    .B1(_02228_),
    .B2(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_2 _18162_ (.A(_02736_),
    .X(_03450_));
 sky130_fd_sc_hd__buf_2 _18163_ (.A(_02740_),
    .X(_03451_));
 sky130_fd_sc_hd__a22oi_4 _18164_ (.A1(\CPU_Xreg_value_a4[23][18] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][18] ),
    .B2(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__inv_2 _18165_ (.A(\CPU_Xreg_value_a4[19][18] ),
    .Y(_03453_));
 sky130_fd_sc_hd__buf_2 _18166_ (.A(_02744_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_2 _18167_ (.A(_02747_),
    .X(_03455_));
 sky130_fd_sc_hd__o22a_4 _18168_ (.A1(_03453_),
    .A2(_03454_),
    .B1(_02252_),
    .B2(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__and4_4 _18169_ (.A(_03446_),
    .B(_03449_),
    .C(_03452_),
    .D(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_2 _18170_ (.A(_02752_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_2 _18171_ (.A(_02756_),
    .X(_03459_));
 sky130_fd_sc_hd__o22a_4 _18172_ (.A1(_02218_),
    .A2(_03458_),
    .B1(_02250_),
    .B2(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__inv_2 _18173_ (.A(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__inv_2 _18174_ (.A(\CPU_Xreg_value_a4[25][18] ),
    .Y(_03462_));
 sky130_fd_sc_hd__buf_2 _18175_ (.A(_02761_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_2 _18176_ (.A(_02765_),
    .X(_03464_));
 sky130_fd_sc_hd__a2bb2o_4 _18177_ (.A1_N(_03462_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][18] ),
    .B2(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__buf_2 _18178_ (.A(_02771_),
    .X(_03466_));
 sky130_fd_sc_hd__inv_2 _18179_ (.A(\CPU_Xreg_value_a4[17][18] ),
    .Y(_03467_));
 sky130_fd_sc_hd__buf_2 _18180_ (.A(_02778_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_2 _18181_ (.A(_02783_),
    .X(_03469_));
 sky130_fd_sc_hd__a2bb2o_4 _18182_ (.A1_N(_03467_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][18] ),
    .B2(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__a211o_4 _18183_ (.A1(\CPU_Xreg_value_a4[13][18] ),
    .A2(_03466_),
    .B1(_03379_),
    .C1(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__inv_2 _18184_ (.A(\CPU_Xreg_value_a4[18][18] ),
    .Y(_03472_));
 sky130_fd_sc_hd__buf_2 _18185_ (.A(_02789_),
    .X(_03473_));
 sky130_fd_sc_hd__buf_2 _18186_ (.A(_02793_),
    .X(_03474_));
 sky130_fd_sc_hd__a2bb2o_4 _18187_ (.A1_N(_03472_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][18] ),
    .B2(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__buf_2 _18188_ (.A(_02797_),
    .X(_03476_));
 sky130_fd_sc_hd__buf_2 _18189_ (.A(_02800_),
    .X(_03477_));
 sky130_fd_sc_hd__o22a_4 _18190_ (.A1(_02226_),
    .A2(_03476_),
    .B1(_02235_),
    .B2(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__inv_2 _18191_ (.A(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__inv_2 _18192_ (.A(\CPU_Xreg_value_a4[21][18] ),
    .Y(_03480_));
 sky130_fd_sc_hd__buf_2 _18193_ (.A(_02805_),
    .X(_03481_));
 sky130_fd_sc_hd__buf_2 _18194_ (.A(_02809_),
    .X(_03482_));
 sky130_fd_sc_hd__a2bb2o_4 _18195_ (.A1_N(_03480_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][18] ),
    .B2(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__inv_2 _18196_ (.A(\CPU_Xreg_value_a4[27][18] ),
    .Y(_03484_));
 sky130_fd_sc_hd__buf_2 _18197_ (.A(_02813_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_2 _18198_ (.A(_02817_),
    .X(_03486_));
 sky130_fd_sc_hd__a2bb2o_4 _18199_ (.A1_N(_03484_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][18] ),
    .B2(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__or4_4 _18200_ (.A(_03475_),
    .B(_03479_),
    .C(_03483_),
    .D(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__or4_4 _18201_ (.A(_03461_),
    .B(_03465_),
    .C(_03471_),
    .D(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__inv_2 _18202_ (.A(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__buf_2 _18203_ (.A(_02823_),
    .X(_03491_));
 sky130_fd_sc_hd__a32o_4 _18204_ (.A1(_03442_),
    .A2(_03457_),
    .A3(_03490_),
    .B1(_06121_),
    .B2(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__inv_2 _18205_ (.A(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__o22a_4 _18206_ (.A1(_06680_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03493_),
    .X(\CPU_src2_value_a2[18] ));
 sky130_fd_sc_hd__o22a_4 _18207_ (.A1(_02271_),
    .A2(_03430_),
    .B1(_02282_),
    .B2(_03431_),
    .X(_03494_));
 sky130_fd_sc_hd__a22oi_4 _18208_ (.A1(\CPU_Xreg_value_a4[16][19] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][19] ),
    .B2(_03434_),
    .Y(_03495_));
 sky130_fd_sc_hd__o22a_4 _18209_ (.A1(_02278_),
    .A2(_03436_),
    .B1(_02263_),
    .B2(_03437_),
    .X(_03496_));
 sky130_fd_sc_hd__o22a_4 _18210_ (.A1(_02276_),
    .A2(_03439_),
    .B1(_02279_),
    .B2(_03440_),
    .X(_03497_));
 sky130_fd_sc_hd__and4_4 _18211_ (.A(_03494_),
    .B(_03495_),
    .C(_03496_),
    .D(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__inv_2 _18212_ (.A(\CPU_Xreg_value_a4[26][19] ),
    .Y(_03499_));
 sky130_fd_sc_hd__o22a_4 _18213_ (.A1(_03499_),
    .A2(_03444_),
    .B1(_02264_),
    .B2(_03445_),
    .X(_03500_));
 sky130_fd_sc_hd__o22a_4 _18214_ (.A1(_02281_),
    .A2(_03447_),
    .B1(_02270_),
    .B2(_03448_),
    .X(_03501_));
 sky130_fd_sc_hd__a22oi_4 _18215_ (.A1(\CPU_Xreg_value_a4[23][19] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][19] ),
    .B2(_03451_),
    .Y(_03502_));
 sky130_fd_sc_hd__inv_2 _18216_ (.A(\CPU_Xreg_value_a4[19][19] ),
    .Y(_03503_));
 sky130_fd_sc_hd__o22a_4 _18217_ (.A1(_03503_),
    .A2(_03454_),
    .B1(_02285_),
    .B2(_03455_),
    .X(_03504_));
 sky130_fd_sc_hd__and4_4 _18218_ (.A(_03500_),
    .B(_03501_),
    .C(_03502_),
    .D(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__o22a_4 _18219_ (.A1(_02259_),
    .A2(_03458_),
    .B1(_02284_),
    .B2(_03459_),
    .X(_03506_));
 sky130_fd_sc_hd__inv_2 _18220_ (.A(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__inv_2 _18221_ (.A(\CPU_Xreg_value_a4[25][19] ),
    .Y(_03508_));
 sky130_fd_sc_hd__a2bb2o_4 _18222_ (.A1_N(_03508_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][19] ),
    .B2(_03464_),
    .X(_03509_));
 sky130_fd_sc_hd__inv_2 _18223_ (.A(\CPU_Xreg_value_a4[17][19] ),
    .Y(_03510_));
 sky130_fd_sc_hd__a2bb2o_4 _18224_ (.A1_N(_03510_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][19] ),
    .B2(_03469_),
    .X(_03511_));
 sky130_fd_sc_hd__a211o_4 _18225_ (.A1(\CPU_Xreg_value_a4[13][19] ),
    .A2(_03466_),
    .B1(_03379_),
    .C1(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__inv_2 _18226_ (.A(\CPU_Xreg_value_a4[18][19] ),
    .Y(_03513_));
 sky130_fd_sc_hd__a2bb2o_4 _18227_ (.A1_N(_03513_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][19] ),
    .B2(_03474_),
    .X(_03514_));
 sky130_fd_sc_hd__o22a_4 _18228_ (.A1(_02267_),
    .A2(_03476_),
    .B1(_02275_),
    .B2(_03477_),
    .X(_03515_));
 sky130_fd_sc_hd__inv_2 _18229_ (.A(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _18230_ (.A(\CPU_Xreg_value_a4[21][19] ),
    .Y(_03517_));
 sky130_fd_sc_hd__a2bb2o_4 _18231_ (.A1_N(_03517_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][19] ),
    .B2(_03482_),
    .X(_03518_));
 sky130_fd_sc_hd__inv_2 _18232_ (.A(\CPU_Xreg_value_a4[27][19] ),
    .Y(_03519_));
 sky130_fd_sc_hd__a2bb2o_4 _18233_ (.A1_N(_03519_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][19] ),
    .B2(_03486_),
    .X(_03520_));
 sky130_fd_sc_hd__or4_4 _18234_ (.A(_03514_),
    .B(_03516_),
    .C(_03518_),
    .D(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__or4_4 _18235_ (.A(_03507_),
    .B(_03509_),
    .C(_03512_),
    .D(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__inv_2 _18236_ (.A(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__a32o_4 _18237_ (.A1(_03498_),
    .A2(_03505_),
    .A3(_03523_),
    .B1(_06120_),
    .B2(_03491_),
    .X(_03524_));
 sky130_fd_sc_hd__inv_2 _18238_ (.A(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__o22a_4 _18239_ (.A1(_06671_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03525_),
    .X(\CPU_src2_value_a2[19] ));
 sky130_fd_sc_hd__o22a_4 _18240_ (.A1(_02299_),
    .A2(_03430_),
    .B1(_02310_),
    .B2(_03431_),
    .X(_03526_));
 sky130_fd_sc_hd__a22oi_4 _18241_ (.A1(\CPU_Xreg_value_a4[16][20] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][20] ),
    .B2(_03434_),
    .Y(_03527_));
 sky130_fd_sc_hd__o22a_4 _18242_ (.A1(_02306_),
    .A2(_03436_),
    .B1(_02292_),
    .B2(_03437_),
    .X(_03528_));
 sky130_fd_sc_hd__o22a_4 _18243_ (.A1(_02304_),
    .A2(_03439_),
    .B1(_02307_),
    .B2(_03440_),
    .X(_03529_));
 sky130_fd_sc_hd__and4_4 _18244_ (.A(_03526_),
    .B(_03527_),
    .C(_03528_),
    .D(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__inv_2 _18245_ (.A(\CPU_Xreg_value_a4[26][20] ),
    .Y(_03531_));
 sky130_fd_sc_hd__o22a_4 _18246_ (.A1(_03531_),
    .A2(_03444_),
    .B1(_02293_),
    .B2(_03445_),
    .X(_03532_));
 sky130_fd_sc_hd__o22a_4 _18247_ (.A1(_02309_),
    .A2(_03447_),
    .B1(_02298_),
    .B2(_03448_),
    .X(_03533_));
 sky130_fd_sc_hd__a22oi_4 _18248_ (.A1(\CPU_Xreg_value_a4[23][20] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][20] ),
    .B2(_03451_),
    .Y(_03534_));
 sky130_fd_sc_hd__inv_2 _18249_ (.A(\CPU_Xreg_value_a4[19][20] ),
    .Y(_03535_));
 sky130_fd_sc_hd__o22a_4 _18250_ (.A1(_03535_),
    .A2(_03454_),
    .B1(_02313_),
    .B2(_03455_),
    .X(_03536_));
 sky130_fd_sc_hd__and4_4 _18251_ (.A(_03532_),
    .B(_03533_),
    .C(_03534_),
    .D(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__o22a_4 _18252_ (.A1(_02290_),
    .A2(_03458_),
    .B1(_02312_),
    .B2(_03459_),
    .X(_03538_));
 sky130_fd_sc_hd__inv_2 _18253_ (.A(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__inv_2 _18254_ (.A(\CPU_Xreg_value_a4[25][20] ),
    .Y(_03540_));
 sky130_fd_sc_hd__a2bb2o_4 _18255_ (.A1_N(_03540_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][20] ),
    .B2(_03464_),
    .X(_03541_));
 sky130_fd_sc_hd__inv_2 _18256_ (.A(\CPU_Xreg_value_a4[17][20] ),
    .Y(_03542_));
 sky130_fd_sc_hd__a2bb2o_4 _18257_ (.A1_N(_03542_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][20] ),
    .B2(_03469_),
    .X(_03543_));
 sky130_fd_sc_hd__a211o_4 _18258_ (.A1(\CPU_Xreg_value_a4[13][20] ),
    .A2(_03466_),
    .B1(_03379_),
    .C1(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__inv_2 _18259_ (.A(\CPU_Xreg_value_a4[18][20] ),
    .Y(_03545_));
 sky130_fd_sc_hd__a2bb2o_4 _18260_ (.A1_N(_03545_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][20] ),
    .B2(_03474_),
    .X(_03546_));
 sky130_fd_sc_hd__o22a_4 _18261_ (.A1(_02296_),
    .A2(_03476_),
    .B1(_02303_),
    .B2(_03477_),
    .X(_03547_));
 sky130_fd_sc_hd__inv_2 _18262_ (.A(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__inv_2 _18263_ (.A(\CPU_Xreg_value_a4[21][20] ),
    .Y(_03549_));
 sky130_fd_sc_hd__a2bb2o_4 _18264_ (.A1_N(_03549_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][20] ),
    .B2(_03482_),
    .X(_03550_));
 sky130_fd_sc_hd__inv_2 _18265_ (.A(\CPU_Xreg_value_a4[27][20] ),
    .Y(_03551_));
 sky130_fd_sc_hd__a2bb2o_4 _18266_ (.A1_N(_03551_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][20] ),
    .B2(_03486_),
    .X(_03552_));
 sky130_fd_sc_hd__or4_4 _18267_ (.A(_03546_),
    .B(_03548_),
    .C(_03550_),
    .D(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__or4_4 _18268_ (.A(_03539_),
    .B(_03541_),
    .C(_03544_),
    .D(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__inv_2 _18269_ (.A(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__a32o_4 _18270_ (.A1(_03530_),
    .A2(_03537_),
    .A3(_03555_),
    .B1(_06117_),
    .B2(_03491_),
    .X(_03556_));
 sky130_fd_sc_hd__inv_2 _18271_ (.A(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__o22a_4 _18272_ (.A1(_06649_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03557_),
    .X(\CPU_src2_value_a2[20] ));
 sky130_fd_sc_hd__o22a_4 _18273_ (.A1(_02327_),
    .A2(_03430_),
    .B1(_02338_),
    .B2(_03431_),
    .X(_03558_));
 sky130_fd_sc_hd__a22oi_4 _18274_ (.A1(\CPU_Xreg_value_a4[16][21] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][21] ),
    .B2(_03434_),
    .Y(_03559_));
 sky130_fd_sc_hd__o22a_4 _18275_ (.A1(_02334_),
    .A2(_03436_),
    .B1(_02320_),
    .B2(_03437_),
    .X(_03560_));
 sky130_fd_sc_hd__o22a_4 _18276_ (.A1(_02332_),
    .A2(_03439_),
    .B1(_02335_),
    .B2(_03440_),
    .X(_03561_));
 sky130_fd_sc_hd__and4_4 _18277_ (.A(_03558_),
    .B(_03559_),
    .C(_03560_),
    .D(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__inv_2 _18278_ (.A(\CPU_Xreg_value_a4[26][21] ),
    .Y(_03563_));
 sky130_fd_sc_hd__o22a_4 _18279_ (.A1(_03563_),
    .A2(_03444_),
    .B1(_02321_),
    .B2(_03445_),
    .X(_03564_));
 sky130_fd_sc_hd__o22a_4 _18280_ (.A1(_02337_),
    .A2(_03447_),
    .B1(_02326_),
    .B2(_03448_),
    .X(_03565_));
 sky130_fd_sc_hd__a22oi_4 _18281_ (.A1(\CPU_Xreg_value_a4[23][21] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][21] ),
    .B2(_03451_),
    .Y(_03566_));
 sky130_fd_sc_hd__inv_2 _18282_ (.A(\CPU_Xreg_value_a4[19][21] ),
    .Y(_03567_));
 sky130_fd_sc_hd__o22a_4 _18283_ (.A1(_03567_),
    .A2(_03454_),
    .B1(_02341_),
    .B2(_03455_),
    .X(_03568_));
 sky130_fd_sc_hd__and4_4 _18284_ (.A(_03564_),
    .B(_03565_),
    .C(_03566_),
    .D(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__o22a_4 _18285_ (.A1(_02318_),
    .A2(_03458_),
    .B1(_02340_),
    .B2(_03459_),
    .X(_03570_));
 sky130_fd_sc_hd__inv_2 _18286_ (.A(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__inv_2 _18287_ (.A(\CPU_Xreg_value_a4[25][21] ),
    .Y(_03572_));
 sky130_fd_sc_hd__a2bb2o_4 _18288_ (.A1_N(_03572_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][21] ),
    .B2(_03464_),
    .X(_03573_));
 sky130_fd_sc_hd__inv_2 _18289_ (.A(\CPU_Xreg_value_a4[17][21] ),
    .Y(_03574_));
 sky130_fd_sc_hd__a2bb2o_4 _18290_ (.A1_N(_03574_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][21] ),
    .B2(_03469_),
    .X(_03575_));
 sky130_fd_sc_hd__a211o_4 _18291_ (.A1(\CPU_Xreg_value_a4[13][21] ),
    .A2(_03466_),
    .B1(_03379_),
    .C1(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__inv_2 _18292_ (.A(\CPU_Xreg_value_a4[18][21] ),
    .Y(_03577_));
 sky130_fd_sc_hd__a2bb2o_4 _18293_ (.A1_N(_03577_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][21] ),
    .B2(_03474_),
    .X(_03578_));
 sky130_fd_sc_hd__o22a_4 _18294_ (.A1(_02324_),
    .A2(_03476_),
    .B1(_02331_),
    .B2(_03477_),
    .X(_03579_));
 sky130_fd_sc_hd__inv_2 _18295_ (.A(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__inv_2 _18296_ (.A(\CPU_Xreg_value_a4[21][21] ),
    .Y(_03581_));
 sky130_fd_sc_hd__a2bb2o_4 _18297_ (.A1_N(_03581_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][21] ),
    .B2(_03482_),
    .X(_03582_));
 sky130_fd_sc_hd__inv_2 _18298_ (.A(\CPU_Xreg_value_a4[27][21] ),
    .Y(_03583_));
 sky130_fd_sc_hd__a2bb2o_4 _18299_ (.A1_N(_03583_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][21] ),
    .B2(_03486_),
    .X(_03584_));
 sky130_fd_sc_hd__or4_4 _18300_ (.A(_03578_),
    .B(_03580_),
    .C(_03582_),
    .D(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__or4_4 _18301_ (.A(_03571_),
    .B(_03573_),
    .C(_03576_),
    .D(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__inv_2 _18302_ (.A(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__a32o_4 _18303_ (.A1(_03562_),
    .A2(_03569_),
    .A3(_03587_),
    .B1(_06116_),
    .B2(_03491_),
    .X(_03588_));
 sky130_fd_sc_hd__inv_2 _18304_ (.A(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__o22a_4 _18305_ (.A1(_06640_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03589_),
    .X(\CPU_src2_value_a2[21] ));
 sky130_fd_sc_hd__o22a_4 _18306_ (.A1(_02355_),
    .A2(_03430_),
    .B1(_02366_),
    .B2(_03431_),
    .X(_03590_));
 sky130_fd_sc_hd__a22oi_4 _18307_ (.A1(\CPU_Xreg_value_a4[16][22] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][22] ),
    .B2(_03434_),
    .Y(_03591_));
 sky130_fd_sc_hd__o22a_4 _18308_ (.A1(_02362_),
    .A2(_03436_),
    .B1(_02348_),
    .B2(_03437_),
    .X(_03592_));
 sky130_fd_sc_hd__o22a_4 _18309_ (.A1(_02360_),
    .A2(_03439_),
    .B1(_02363_),
    .B2(_03440_),
    .X(_03593_));
 sky130_fd_sc_hd__and4_4 _18310_ (.A(_03590_),
    .B(_03591_),
    .C(_03592_),
    .D(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__inv_2 _18311_ (.A(\CPU_Xreg_value_a4[26][22] ),
    .Y(_03595_));
 sky130_fd_sc_hd__o22a_4 _18312_ (.A1(_03595_),
    .A2(_03444_),
    .B1(_02349_),
    .B2(_03445_),
    .X(_03596_));
 sky130_fd_sc_hd__o22a_4 _18313_ (.A1(_02365_),
    .A2(_03447_),
    .B1(_02354_),
    .B2(_03448_),
    .X(_03597_));
 sky130_fd_sc_hd__a22oi_4 _18314_ (.A1(\CPU_Xreg_value_a4[23][22] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][22] ),
    .B2(_03451_),
    .Y(_03598_));
 sky130_fd_sc_hd__inv_2 _18315_ (.A(\CPU_Xreg_value_a4[19][22] ),
    .Y(_03599_));
 sky130_fd_sc_hd__o22a_4 _18316_ (.A1(_03599_),
    .A2(_03454_),
    .B1(_02369_),
    .B2(_03455_),
    .X(_03600_));
 sky130_fd_sc_hd__and4_4 _18317_ (.A(_03596_),
    .B(_03597_),
    .C(_03598_),
    .D(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__o22a_4 _18318_ (.A1(_02346_),
    .A2(_03458_),
    .B1(_02368_),
    .B2(_03459_),
    .X(_03602_));
 sky130_fd_sc_hd__inv_2 _18319_ (.A(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__inv_2 _18320_ (.A(\CPU_Xreg_value_a4[25][22] ),
    .Y(_03604_));
 sky130_fd_sc_hd__a2bb2o_4 _18321_ (.A1_N(_03604_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][22] ),
    .B2(_03464_),
    .X(_03605_));
 sky130_fd_sc_hd__buf_2 _18322_ (.A(_02774_),
    .X(_03606_));
 sky130_fd_sc_hd__inv_2 _18323_ (.A(\CPU_Xreg_value_a4[17][22] ),
    .Y(_03607_));
 sky130_fd_sc_hd__a2bb2o_4 _18324_ (.A1_N(_03607_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][22] ),
    .B2(_03469_),
    .X(_03608_));
 sky130_fd_sc_hd__a211o_4 _18325_ (.A1(\CPU_Xreg_value_a4[13][22] ),
    .A2(_03466_),
    .B1(_03606_),
    .C1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__inv_2 _18326_ (.A(\CPU_Xreg_value_a4[18][22] ),
    .Y(_03610_));
 sky130_fd_sc_hd__a2bb2o_4 _18327_ (.A1_N(_03610_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][22] ),
    .B2(_03474_),
    .X(_03611_));
 sky130_fd_sc_hd__o22a_4 _18328_ (.A1(_02352_),
    .A2(_03476_),
    .B1(_02359_),
    .B2(_03477_),
    .X(_03612_));
 sky130_fd_sc_hd__inv_2 _18329_ (.A(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__inv_2 _18330_ (.A(\CPU_Xreg_value_a4[21][22] ),
    .Y(_03614_));
 sky130_fd_sc_hd__a2bb2o_4 _18331_ (.A1_N(_03614_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][22] ),
    .B2(_03482_),
    .X(_03615_));
 sky130_fd_sc_hd__inv_2 _18332_ (.A(\CPU_Xreg_value_a4[27][22] ),
    .Y(_03616_));
 sky130_fd_sc_hd__a2bb2o_4 _18333_ (.A1_N(_03616_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][22] ),
    .B2(_03486_),
    .X(_03617_));
 sky130_fd_sc_hd__or4_4 _18334_ (.A(_03611_),
    .B(_03613_),
    .C(_03615_),
    .D(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__or4_4 _18335_ (.A(_03603_),
    .B(_03605_),
    .C(_03609_),
    .D(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__inv_2 _18336_ (.A(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__a32o_4 _18337_ (.A1(_03594_),
    .A2(_03601_),
    .A3(_03620_),
    .B1(_06115_),
    .B2(_03491_),
    .X(_03621_));
 sky130_fd_sc_hd__inv_2 _18338_ (.A(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__o22a_4 _18339_ (.A1(_06625_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03622_),
    .X(\CPU_src2_value_a2[22] ));
 sky130_fd_sc_hd__o22a_4 _18340_ (.A1(_02384_),
    .A2(_03430_),
    .B1(_02395_),
    .B2(_03431_),
    .X(_03623_));
 sky130_fd_sc_hd__a22oi_4 _18341_ (.A1(\CPU_Xreg_value_a4[16][23] ),
    .A2(_03433_),
    .B1(\CPU_Xreg_value_a4[30][23] ),
    .B2(_03434_),
    .Y(_03624_));
 sky130_fd_sc_hd__o22a_4 _18342_ (.A1(_02391_),
    .A2(_03436_),
    .B1(_02376_),
    .B2(_03437_),
    .X(_03625_));
 sky130_fd_sc_hd__o22a_4 _18343_ (.A1(_02389_),
    .A2(_03439_),
    .B1(_02392_),
    .B2(_03440_),
    .X(_03626_));
 sky130_fd_sc_hd__and4_4 _18344_ (.A(_03623_),
    .B(_03624_),
    .C(_03625_),
    .D(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__inv_2 _18345_ (.A(\CPU_Xreg_value_a4[26][23] ),
    .Y(_03628_));
 sky130_fd_sc_hd__o22a_4 _18346_ (.A1(_03628_),
    .A2(_03444_),
    .B1(_02377_),
    .B2(_03445_),
    .X(_03629_));
 sky130_fd_sc_hd__o22a_4 _18347_ (.A1(_02394_),
    .A2(_03447_),
    .B1(_02383_),
    .B2(_03448_),
    .X(_03630_));
 sky130_fd_sc_hd__a22oi_4 _18348_ (.A1(\CPU_Xreg_value_a4[23][23] ),
    .A2(_03450_),
    .B1(\CPU_Xreg_value_a4[31][23] ),
    .B2(_03451_),
    .Y(_03631_));
 sky130_fd_sc_hd__inv_2 _18349_ (.A(\CPU_Xreg_value_a4[19][23] ),
    .Y(_03632_));
 sky130_fd_sc_hd__o22a_4 _18350_ (.A1(_03632_),
    .A2(_03454_),
    .B1(_02398_),
    .B2(_03455_),
    .X(_03633_));
 sky130_fd_sc_hd__and4_4 _18351_ (.A(_03629_),
    .B(_03630_),
    .C(_03631_),
    .D(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o22a_4 _18352_ (.A1(_02374_),
    .A2(_03458_),
    .B1(_02397_),
    .B2(_03459_),
    .X(_03635_));
 sky130_fd_sc_hd__inv_2 _18353_ (.A(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__inv_2 _18354_ (.A(\CPU_Xreg_value_a4[25][23] ),
    .Y(_03637_));
 sky130_fd_sc_hd__a2bb2o_4 _18355_ (.A1_N(_03637_),
    .A2_N(_03463_),
    .B1(\CPU_Xreg_value_a4[24][23] ),
    .B2(_03464_),
    .X(_03638_));
 sky130_fd_sc_hd__inv_2 _18356_ (.A(\CPU_Xreg_value_a4[17][23] ),
    .Y(_03639_));
 sky130_fd_sc_hd__a2bb2o_4 _18357_ (.A1_N(_03639_),
    .A2_N(_03468_),
    .B1(\CPU_Xreg_value_a4[22][23] ),
    .B2(_03469_),
    .X(_03640_));
 sky130_fd_sc_hd__a211o_4 _18358_ (.A1(\CPU_Xreg_value_a4[13][23] ),
    .A2(_03466_),
    .B1(_03606_),
    .C1(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__inv_2 _18359_ (.A(\CPU_Xreg_value_a4[18][23] ),
    .Y(_03642_));
 sky130_fd_sc_hd__a2bb2o_4 _18360_ (.A1_N(_03642_),
    .A2_N(_03473_),
    .B1(\CPU_Xreg_value_a4[28][23] ),
    .B2(_03474_),
    .X(_03643_));
 sky130_fd_sc_hd__o22a_4 _18361_ (.A1(_02380_),
    .A2(_03476_),
    .B1(_02388_),
    .B2(_03477_),
    .X(_03644_));
 sky130_fd_sc_hd__inv_2 _18362_ (.A(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__inv_2 _18363_ (.A(\CPU_Xreg_value_a4[21][23] ),
    .Y(_03646_));
 sky130_fd_sc_hd__a2bb2o_4 _18364_ (.A1_N(_03646_),
    .A2_N(_03481_),
    .B1(\CPU_Xreg_value_a4[20][23] ),
    .B2(_03482_),
    .X(_03647_));
 sky130_fd_sc_hd__inv_2 _18365_ (.A(\CPU_Xreg_value_a4[27][23] ),
    .Y(_03648_));
 sky130_fd_sc_hd__a2bb2o_4 _18366_ (.A1_N(_03648_),
    .A2_N(_03485_),
    .B1(\CPU_Xreg_value_a4[29][23] ),
    .B2(_03486_),
    .X(_03649_));
 sky130_fd_sc_hd__or4_4 _18367_ (.A(_03643_),
    .B(_03645_),
    .C(_03647_),
    .D(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__or4_4 _18368_ (.A(_03636_),
    .B(_03638_),
    .C(_03641_),
    .D(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__inv_2 _18369_ (.A(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a32o_4 _18370_ (.A1(_03627_),
    .A2(_03634_),
    .A3(_03652_),
    .B1(_06114_),
    .B2(_03491_),
    .X(_03653_));
 sky130_fd_sc_hd__inv_2 _18371_ (.A(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__o22a_4 _18372_ (.A1(_06617_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03654_),
    .X(\CPU_src2_value_a2[23] ));
 sky130_fd_sc_hd__buf_2 _18373_ (.A(_02668_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_2 _18374_ (.A(_02671_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_2 _18375_ (.A(_02680_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_2 _18376_ (.A(_02685_),
    .X(_03658_));
 sky130_fd_sc_hd__o22a_4 _18377_ (.A1(_02417_),
    .A2(_03657_),
    .B1(_02434_),
    .B2(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_2 _18378_ (.A(_02692_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_2 _18379_ (.A(_02698_),
    .X(_03661_));
 sky130_fd_sc_hd__a22oi_4 _18380_ (.A1(\CPU_Xreg_value_a4[16][24] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][24] ),
    .B2(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__buf_2 _18381_ (.A(_02703_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_2 _18382_ (.A(_02707_),
    .X(_03664_));
 sky130_fd_sc_hd__o22a_4 _18383_ (.A1(_02427_),
    .A2(_03663_),
    .B1(_02407_),
    .B2(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__buf_2 _18384_ (.A(_02711_),
    .X(_03666_));
 sky130_fd_sc_hd__buf_2 _18385_ (.A(_02714_),
    .X(_03667_));
 sky130_fd_sc_hd__o22a_4 _18386_ (.A1(_02424_),
    .A2(_03666_),
    .B1(_02429_),
    .B2(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__and4_4 _18387_ (.A(_03659_),
    .B(_03662_),
    .C(_03665_),
    .D(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__inv_2 _18388_ (.A(\CPU_Xreg_value_a4[26][24] ),
    .Y(_03670_));
 sky130_fd_sc_hd__buf_2 _18389_ (.A(_02720_),
    .X(_03671_));
 sky130_fd_sc_hd__buf_2 _18390_ (.A(_02723_),
    .X(_03672_));
 sky130_fd_sc_hd__o22a_4 _18391_ (.A1(_03670_),
    .A2(_03671_),
    .B1(_02409_),
    .B2(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__buf_2 _18392_ (.A(_02727_),
    .X(_03674_));
 sky130_fd_sc_hd__buf_2 _18393_ (.A(_02730_),
    .X(_03675_));
 sky130_fd_sc_hd__o22a_4 _18394_ (.A1(_02432_),
    .A2(_03674_),
    .B1(_02415_),
    .B2(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__buf_2 _18395_ (.A(_02735_),
    .X(_03677_));
 sky130_fd_sc_hd__buf_2 _18396_ (.A(_02739_),
    .X(_03678_));
 sky130_fd_sc_hd__a22oi_4 _18397_ (.A1(\CPU_Xreg_value_a4[23][24] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][24] ),
    .B2(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__inv_2 _18398_ (.A(\CPU_Xreg_value_a4[19][24] ),
    .Y(_03680_));
 sky130_fd_sc_hd__buf_2 _18399_ (.A(_02743_),
    .X(_03681_));
 sky130_fd_sc_hd__buf_2 _18400_ (.A(_02746_),
    .X(_03682_));
 sky130_fd_sc_hd__o22a_4 _18401_ (.A1(_03680_),
    .A2(_03681_),
    .B1(_02439_),
    .B2(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__and4_4 _18402_ (.A(_03673_),
    .B(_03676_),
    .C(_03679_),
    .D(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_2 _18403_ (.A(_02751_),
    .X(_03685_));
 sky130_fd_sc_hd__buf_2 _18404_ (.A(_02755_),
    .X(_03686_));
 sky130_fd_sc_hd__o22a_4 _18405_ (.A1(_02405_),
    .A2(_03685_),
    .B1(_02437_),
    .B2(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__inv_2 _18406_ (.A(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__inv_2 _18407_ (.A(\CPU_Xreg_value_a4[25][24] ),
    .Y(_03689_));
 sky130_fd_sc_hd__buf_2 _18408_ (.A(_02760_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_2 _18409_ (.A(_02764_),
    .X(_03691_));
 sky130_fd_sc_hd__a2bb2o_4 _18410_ (.A1_N(_03689_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][24] ),
    .B2(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_2 _18411_ (.A(_02770_),
    .X(_03693_));
 sky130_fd_sc_hd__inv_2 _18412_ (.A(\CPU_Xreg_value_a4[17][24] ),
    .Y(_03694_));
 sky130_fd_sc_hd__buf_2 _18413_ (.A(_02777_),
    .X(_03695_));
 sky130_fd_sc_hd__buf_2 _18414_ (.A(_02782_),
    .X(_03696_));
 sky130_fd_sc_hd__a2bb2o_4 _18415_ (.A1_N(_03694_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][24] ),
    .B2(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__a211o_4 _18416_ (.A1(\CPU_Xreg_value_a4[13][24] ),
    .A2(_03693_),
    .B1(_03606_),
    .C1(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__inv_2 _18417_ (.A(\CPU_Xreg_value_a4[18][24] ),
    .Y(_03699_));
 sky130_fd_sc_hd__buf_2 _18418_ (.A(_02788_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_2 _18419_ (.A(_02792_),
    .X(_03701_));
 sky130_fd_sc_hd__a2bb2o_4 _18420_ (.A1_N(_03699_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][24] ),
    .B2(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_2 _18421_ (.A(_02796_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_2 _18422_ (.A(_02799_),
    .X(_03704_));
 sky130_fd_sc_hd__o22a_4 _18423_ (.A1(_02413_),
    .A2(_03703_),
    .B1(_02422_),
    .B2(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__inv_2 _18424_ (.A(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__inv_2 _18425_ (.A(\CPU_Xreg_value_a4[21][24] ),
    .Y(_03707_));
 sky130_fd_sc_hd__buf_2 _18426_ (.A(_02804_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_2 _18427_ (.A(_02808_),
    .X(_03709_));
 sky130_fd_sc_hd__a2bb2o_4 _18428_ (.A1_N(_03707_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][24] ),
    .B2(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__inv_2 _18429_ (.A(\CPU_Xreg_value_a4[27][24] ),
    .Y(_03711_));
 sky130_fd_sc_hd__buf_2 _18430_ (.A(_02812_),
    .X(_03712_));
 sky130_fd_sc_hd__buf_2 _18431_ (.A(_02816_),
    .X(_03713_));
 sky130_fd_sc_hd__a2bb2o_4 _18432_ (.A1_N(_03711_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][24] ),
    .B2(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__or4_4 _18433_ (.A(_03702_),
    .B(_03706_),
    .C(_03710_),
    .D(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__or4_4 _18434_ (.A(_03688_),
    .B(_03692_),
    .C(_03698_),
    .D(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__inv_2 _18435_ (.A(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__buf_2 _18436_ (.A(_02775_),
    .X(_03718_));
 sky130_fd_sc_hd__a32o_4 _18437_ (.A1(_03669_),
    .A2(_03684_),
    .A3(_03717_),
    .B1(_06113_),
    .B2(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__inv_2 _18438_ (.A(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__o22a_4 _18439_ (.A1(_06597_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03720_),
    .X(\CPU_src2_value_a2[24] ));
 sky130_fd_sc_hd__o22a_4 _18440_ (.A1(_02458_),
    .A2(_03657_),
    .B1(_02469_),
    .B2(_03658_),
    .X(_03721_));
 sky130_fd_sc_hd__a22oi_4 _18441_ (.A1(\CPU_Xreg_value_a4[16][25] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][25] ),
    .B2(_03661_),
    .Y(_03722_));
 sky130_fd_sc_hd__o22a_4 _18442_ (.A1(_02465_),
    .A2(_03663_),
    .B1(_02450_),
    .B2(_03664_),
    .X(_03723_));
 sky130_fd_sc_hd__o22a_4 _18443_ (.A1(_02463_),
    .A2(_03666_),
    .B1(_02466_),
    .B2(_03667_),
    .X(_03724_));
 sky130_fd_sc_hd__and4_4 _18444_ (.A(_03721_),
    .B(_03722_),
    .C(_03723_),
    .D(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__inv_2 _18445_ (.A(\CPU_Xreg_value_a4[26][25] ),
    .Y(_03726_));
 sky130_fd_sc_hd__o22a_4 _18446_ (.A1(_03726_),
    .A2(_03671_),
    .B1(_02451_),
    .B2(_03672_),
    .X(_03727_));
 sky130_fd_sc_hd__o22a_4 _18447_ (.A1(_02468_),
    .A2(_03674_),
    .B1(_02457_),
    .B2(_03675_),
    .X(_03728_));
 sky130_fd_sc_hd__a22oi_4 _18448_ (.A1(\CPU_Xreg_value_a4[23][25] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][25] ),
    .B2(_03678_),
    .Y(_03729_));
 sky130_fd_sc_hd__inv_2 _18449_ (.A(\CPU_Xreg_value_a4[19][25] ),
    .Y(_03730_));
 sky130_fd_sc_hd__o22a_4 _18450_ (.A1(_03730_),
    .A2(_03681_),
    .B1(_02472_),
    .B2(_03682_),
    .X(_03731_));
 sky130_fd_sc_hd__and4_4 _18451_ (.A(_03727_),
    .B(_03728_),
    .C(_03729_),
    .D(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__o22a_4 _18452_ (.A1(_02446_),
    .A2(_03685_),
    .B1(_02471_),
    .B2(_03686_),
    .X(_03733_));
 sky130_fd_sc_hd__inv_2 _18453_ (.A(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__inv_2 _18454_ (.A(\CPU_Xreg_value_a4[25][25] ),
    .Y(_03735_));
 sky130_fd_sc_hd__a2bb2o_4 _18455_ (.A1_N(_03735_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][25] ),
    .B2(_03691_),
    .X(_03736_));
 sky130_fd_sc_hd__inv_2 _18456_ (.A(\CPU_Xreg_value_a4[17][25] ),
    .Y(_03737_));
 sky130_fd_sc_hd__a2bb2o_4 _18457_ (.A1_N(_03737_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][25] ),
    .B2(_03696_),
    .X(_03738_));
 sky130_fd_sc_hd__a211o_4 _18458_ (.A1(\CPU_Xreg_value_a4[13][25] ),
    .A2(_03693_),
    .B1(_03606_),
    .C1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__inv_2 _18459_ (.A(\CPU_Xreg_value_a4[18][25] ),
    .Y(_03740_));
 sky130_fd_sc_hd__a2bb2o_4 _18460_ (.A1_N(_03740_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][25] ),
    .B2(_03701_),
    .X(_03741_));
 sky130_fd_sc_hd__o22a_4 _18461_ (.A1(_02454_),
    .A2(_03703_),
    .B1(_02462_),
    .B2(_03704_),
    .X(_03742_));
 sky130_fd_sc_hd__inv_2 _18462_ (.A(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__inv_2 _18463_ (.A(\CPU_Xreg_value_a4[21][25] ),
    .Y(_03744_));
 sky130_fd_sc_hd__a2bb2o_4 _18464_ (.A1_N(_03744_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][25] ),
    .B2(_03709_),
    .X(_03745_));
 sky130_fd_sc_hd__inv_2 _18465_ (.A(\CPU_Xreg_value_a4[27][25] ),
    .Y(_03746_));
 sky130_fd_sc_hd__a2bb2o_4 _18466_ (.A1_N(_03746_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][25] ),
    .B2(_03713_),
    .X(_03747_));
 sky130_fd_sc_hd__or4_4 _18467_ (.A(_03741_),
    .B(_03743_),
    .C(_03745_),
    .D(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__or4_4 _18468_ (.A(_03734_),
    .B(_03736_),
    .C(_03739_),
    .D(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__inv_2 _18469_ (.A(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__a32o_4 _18470_ (.A1(_03725_),
    .A2(_03732_),
    .A3(_03750_),
    .B1(_06112_),
    .B2(_03718_),
    .X(_03751_));
 sky130_fd_sc_hd__inv_2 _18471_ (.A(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__o22a_4 _18472_ (.A1(_06587_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03752_),
    .X(\CPU_src2_value_a2[25] ));
 sky130_fd_sc_hd__o22a_4 _18473_ (.A1(_02486_),
    .A2(_03657_),
    .B1(_02497_),
    .B2(_03658_),
    .X(_03753_));
 sky130_fd_sc_hd__a22oi_4 _18474_ (.A1(\CPU_Xreg_value_a4[16][26] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][26] ),
    .B2(_03661_),
    .Y(_03754_));
 sky130_fd_sc_hd__o22a_4 _18475_ (.A1(_02493_),
    .A2(_03663_),
    .B1(_02479_),
    .B2(_03664_),
    .X(_03755_));
 sky130_fd_sc_hd__o22a_4 _18476_ (.A1(_02491_),
    .A2(_03666_),
    .B1(_02494_),
    .B2(_03667_),
    .X(_03756_));
 sky130_fd_sc_hd__and4_4 _18477_ (.A(_03753_),
    .B(_03754_),
    .C(_03755_),
    .D(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__inv_2 _18478_ (.A(\CPU_Xreg_value_a4[26][26] ),
    .Y(_03758_));
 sky130_fd_sc_hd__o22a_4 _18479_ (.A1(_03758_),
    .A2(_03671_),
    .B1(_02480_),
    .B2(_03672_),
    .X(_03759_));
 sky130_fd_sc_hd__o22a_4 _18480_ (.A1(_02496_),
    .A2(_03674_),
    .B1(_02485_),
    .B2(_03675_),
    .X(_03760_));
 sky130_fd_sc_hd__a22oi_4 _18481_ (.A1(\CPU_Xreg_value_a4[23][26] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][26] ),
    .B2(_03678_),
    .Y(_03761_));
 sky130_fd_sc_hd__inv_2 _18482_ (.A(\CPU_Xreg_value_a4[19][26] ),
    .Y(_03762_));
 sky130_fd_sc_hd__o22a_4 _18483_ (.A1(_03762_),
    .A2(_03681_),
    .B1(_02500_),
    .B2(_03682_),
    .X(_03763_));
 sky130_fd_sc_hd__and4_4 _18484_ (.A(_03759_),
    .B(_03760_),
    .C(_03761_),
    .D(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__o22a_4 _18485_ (.A1(_02477_),
    .A2(_03685_),
    .B1(_02499_),
    .B2(_03686_),
    .X(_03765_));
 sky130_fd_sc_hd__inv_2 _18486_ (.A(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__inv_2 _18487_ (.A(\CPU_Xreg_value_a4[25][26] ),
    .Y(_03767_));
 sky130_fd_sc_hd__a2bb2o_4 _18488_ (.A1_N(_03767_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][26] ),
    .B2(_03691_),
    .X(_03768_));
 sky130_fd_sc_hd__inv_2 _18489_ (.A(\CPU_Xreg_value_a4[17][26] ),
    .Y(_03769_));
 sky130_fd_sc_hd__a2bb2o_4 _18490_ (.A1_N(_03769_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][26] ),
    .B2(_03696_),
    .X(_03770_));
 sky130_fd_sc_hd__a211o_4 _18491_ (.A1(\CPU_Xreg_value_a4[13][26] ),
    .A2(_03693_),
    .B1(_03606_),
    .C1(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__inv_2 _18492_ (.A(\CPU_Xreg_value_a4[18][26] ),
    .Y(_03772_));
 sky130_fd_sc_hd__a2bb2o_4 _18493_ (.A1_N(_03772_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][26] ),
    .B2(_03701_),
    .X(_03773_));
 sky130_fd_sc_hd__o22a_4 _18494_ (.A1(_02483_),
    .A2(_03703_),
    .B1(_02490_),
    .B2(_03704_),
    .X(_03774_));
 sky130_fd_sc_hd__inv_2 _18495_ (.A(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__inv_2 _18496_ (.A(\CPU_Xreg_value_a4[21][26] ),
    .Y(_03776_));
 sky130_fd_sc_hd__a2bb2o_4 _18497_ (.A1_N(_03776_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][26] ),
    .B2(_03709_),
    .X(_03777_));
 sky130_fd_sc_hd__inv_2 _18498_ (.A(\CPU_Xreg_value_a4[27][26] ),
    .Y(_03778_));
 sky130_fd_sc_hd__a2bb2o_4 _18499_ (.A1_N(_03778_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][26] ),
    .B2(_03713_),
    .X(_03779_));
 sky130_fd_sc_hd__or4_4 _18500_ (.A(_03773_),
    .B(_03775_),
    .C(_03777_),
    .D(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__or4_4 _18501_ (.A(_03766_),
    .B(_03768_),
    .C(_03771_),
    .D(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__inv_2 _18502_ (.A(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__a32o_4 _18503_ (.A1(_03757_),
    .A2(_03764_),
    .A3(_03782_),
    .B1(_06110_),
    .B2(_03718_),
    .X(_03783_));
 sky130_fd_sc_hd__inv_2 _18504_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__o22a_4 _18505_ (.A1(_06572_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03784_),
    .X(\CPU_src2_value_a2[26] ));
 sky130_fd_sc_hd__o22a_4 _18506_ (.A1(_02514_),
    .A2(_03657_),
    .B1(_02525_),
    .B2(_03658_),
    .X(_03785_));
 sky130_fd_sc_hd__a22oi_4 _18507_ (.A1(\CPU_Xreg_value_a4[16][27] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][27] ),
    .B2(_03661_),
    .Y(_03786_));
 sky130_fd_sc_hd__o22a_4 _18508_ (.A1(_02521_),
    .A2(_03663_),
    .B1(_02507_),
    .B2(_03664_),
    .X(_03787_));
 sky130_fd_sc_hd__o22a_4 _18509_ (.A1(_02519_),
    .A2(_03666_),
    .B1(_02522_),
    .B2(_03667_),
    .X(_03788_));
 sky130_fd_sc_hd__and4_4 _18510_ (.A(_03785_),
    .B(_03786_),
    .C(_03787_),
    .D(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__inv_2 _18511_ (.A(\CPU_Xreg_value_a4[26][27] ),
    .Y(_03790_));
 sky130_fd_sc_hd__o22a_4 _18512_ (.A1(_03790_),
    .A2(_03671_),
    .B1(_02508_),
    .B2(_03672_),
    .X(_03791_));
 sky130_fd_sc_hd__o22a_4 _18513_ (.A1(_02524_),
    .A2(_03674_),
    .B1(_02513_),
    .B2(_03675_),
    .X(_03792_));
 sky130_fd_sc_hd__a22oi_4 _18514_ (.A1(\CPU_Xreg_value_a4[23][27] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][27] ),
    .B2(_03678_),
    .Y(_03793_));
 sky130_fd_sc_hd__inv_2 _18515_ (.A(\CPU_Xreg_value_a4[19][27] ),
    .Y(_03794_));
 sky130_fd_sc_hd__o22a_4 _18516_ (.A1(_03794_),
    .A2(_03681_),
    .B1(_02528_),
    .B2(_03682_),
    .X(_03795_));
 sky130_fd_sc_hd__and4_4 _18517_ (.A(_03791_),
    .B(_03792_),
    .C(_03793_),
    .D(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__o22a_4 _18518_ (.A1(_02505_),
    .A2(_03685_),
    .B1(_02527_),
    .B2(_03686_),
    .X(_03797_));
 sky130_fd_sc_hd__inv_2 _18519_ (.A(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__inv_2 _18520_ (.A(\CPU_Xreg_value_a4[25][27] ),
    .Y(_03799_));
 sky130_fd_sc_hd__a2bb2o_4 _18521_ (.A1_N(_03799_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][27] ),
    .B2(_03691_),
    .X(_03800_));
 sky130_fd_sc_hd__inv_2 _18522_ (.A(\CPU_Xreg_value_a4[17][27] ),
    .Y(_03801_));
 sky130_fd_sc_hd__a2bb2o_4 _18523_ (.A1_N(_03801_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][27] ),
    .B2(_03696_),
    .X(_03802_));
 sky130_fd_sc_hd__a211o_4 _18524_ (.A1(\CPU_Xreg_value_a4[13][27] ),
    .A2(_03693_),
    .B1(_03606_),
    .C1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__inv_2 _18525_ (.A(\CPU_Xreg_value_a4[18][27] ),
    .Y(_03804_));
 sky130_fd_sc_hd__a2bb2o_4 _18526_ (.A1_N(_03804_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][27] ),
    .B2(_03701_),
    .X(_03805_));
 sky130_fd_sc_hd__o22a_4 _18527_ (.A1(_02511_),
    .A2(_03703_),
    .B1(_02518_),
    .B2(_03704_),
    .X(_03806_));
 sky130_fd_sc_hd__inv_2 _18528_ (.A(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__inv_2 _18529_ (.A(\CPU_Xreg_value_a4[21][27] ),
    .Y(_03808_));
 sky130_fd_sc_hd__a2bb2o_4 _18530_ (.A1_N(_03808_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][27] ),
    .B2(_03709_),
    .X(_03809_));
 sky130_fd_sc_hd__inv_2 _18531_ (.A(\CPU_Xreg_value_a4[27][27] ),
    .Y(_03810_));
 sky130_fd_sc_hd__a2bb2o_4 _18532_ (.A1_N(_03810_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][27] ),
    .B2(_03713_),
    .X(_03811_));
 sky130_fd_sc_hd__or4_4 _18533_ (.A(_03805_),
    .B(_03807_),
    .C(_03809_),
    .D(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__or4_4 _18534_ (.A(_03798_),
    .B(_03800_),
    .C(_03803_),
    .D(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__inv_2 _18535_ (.A(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__a32o_4 _18536_ (.A1(_03789_),
    .A2(_03796_),
    .A3(_03814_),
    .B1(_06109_),
    .B2(_03718_),
    .X(_03815_));
 sky130_fd_sc_hd__inv_2 _18537_ (.A(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__o22a_4 _18538_ (.A1(_06562_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03816_),
    .X(\CPU_src2_value_a2[27] ));
 sky130_fd_sc_hd__o22a_4 _18539_ (.A1(_02542_),
    .A2(_03657_),
    .B1(_02553_),
    .B2(_03658_),
    .X(_03817_));
 sky130_fd_sc_hd__a22oi_4 _18540_ (.A1(\CPU_Xreg_value_a4[16][28] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][28] ),
    .B2(_03661_),
    .Y(_03818_));
 sky130_fd_sc_hd__o22a_4 _18541_ (.A1(_02549_),
    .A2(_03663_),
    .B1(_02535_),
    .B2(_03664_),
    .X(_03819_));
 sky130_fd_sc_hd__o22a_4 _18542_ (.A1(_02547_),
    .A2(_03666_),
    .B1(_02550_),
    .B2(_03667_),
    .X(_03820_));
 sky130_fd_sc_hd__and4_4 _18543_ (.A(_03817_),
    .B(_03818_),
    .C(_03819_),
    .D(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__inv_2 _18544_ (.A(\CPU_Xreg_value_a4[26][28] ),
    .Y(_03822_));
 sky130_fd_sc_hd__o22a_4 _18545_ (.A1(_03822_),
    .A2(_03671_),
    .B1(_02536_),
    .B2(_03672_),
    .X(_03823_));
 sky130_fd_sc_hd__o22a_4 _18546_ (.A1(_02552_),
    .A2(_03674_),
    .B1(_02541_),
    .B2(_03675_),
    .X(_03824_));
 sky130_fd_sc_hd__a22oi_4 _18547_ (.A1(\CPU_Xreg_value_a4[23][28] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][28] ),
    .B2(_03678_),
    .Y(_03825_));
 sky130_fd_sc_hd__inv_2 _18548_ (.A(\CPU_Xreg_value_a4[19][28] ),
    .Y(_03826_));
 sky130_fd_sc_hd__o22a_4 _18549_ (.A1(_03826_),
    .A2(_03681_),
    .B1(_02556_),
    .B2(_03682_),
    .X(_03827_));
 sky130_fd_sc_hd__and4_4 _18550_ (.A(_03823_),
    .B(_03824_),
    .C(_03825_),
    .D(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__o22a_4 _18551_ (.A1(_02533_),
    .A2(_03685_),
    .B1(_02555_),
    .B2(_03686_),
    .X(_03829_));
 sky130_fd_sc_hd__inv_2 _18552_ (.A(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__inv_2 _18553_ (.A(\CPU_Xreg_value_a4[25][28] ),
    .Y(_03831_));
 sky130_fd_sc_hd__a2bb2o_4 _18554_ (.A1_N(_03831_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][28] ),
    .B2(_03691_),
    .X(_03832_));
 sky130_fd_sc_hd__inv_2 _18555_ (.A(\CPU_Xreg_value_a4[17][28] ),
    .Y(_03833_));
 sky130_fd_sc_hd__a2bb2o_4 _18556_ (.A1_N(_03833_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][28] ),
    .B2(_03696_),
    .X(_03834_));
 sky130_fd_sc_hd__a211o_4 _18557_ (.A1(\CPU_Xreg_value_a4[13][28] ),
    .A2(_03693_),
    .B1(_02928_),
    .C1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__inv_2 _18558_ (.A(\CPU_Xreg_value_a4[18][28] ),
    .Y(_03836_));
 sky130_fd_sc_hd__a2bb2o_4 _18559_ (.A1_N(_03836_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][28] ),
    .B2(_03701_),
    .X(_03837_));
 sky130_fd_sc_hd__o22a_4 _18560_ (.A1(_02539_),
    .A2(_03703_),
    .B1(_02546_),
    .B2(_03704_),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _18561_ (.A(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__inv_2 _18562_ (.A(\CPU_Xreg_value_a4[21][28] ),
    .Y(_03840_));
 sky130_fd_sc_hd__a2bb2o_4 _18563_ (.A1_N(_03840_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][28] ),
    .B2(_03709_),
    .X(_03841_));
 sky130_fd_sc_hd__inv_2 _18564_ (.A(\CPU_Xreg_value_a4[27][28] ),
    .Y(_03842_));
 sky130_fd_sc_hd__a2bb2o_4 _18565_ (.A1_N(_03842_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][28] ),
    .B2(_03713_),
    .X(_03843_));
 sky130_fd_sc_hd__or4_4 _18566_ (.A(_03837_),
    .B(_03839_),
    .C(_03841_),
    .D(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__or4_4 _18567_ (.A(_03830_),
    .B(_03832_),
    .C(_03835_),
    .D(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__inv_2 _18568_ (.A(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__a32o_4 _18569_ (.A1(_03821_),
    .A2(_03828_),
    .A3(_03846_),
    .B1(_06108_),
    .B2(_03718_),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _18570_ (.A(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__o22a_4 _18571_ (.A1(_06537_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03848_),
    .X(\CPU_src2_value_a2[28] ));
 sky130_fd_sc_hd__o22a_4 _18572_ (.A1(_02570_),
    .A2(_03657_),
    .B1(_02581_),
    .B2(_03658_),
    .X(_03849_));
 sky130_fd_sc_hd__a22oi_4 _18573_ (.A1(\CPU_Xreg_value_a4[16][29] ),
    .A2(_03660_),
    .B1(\CPU_Xreg_value_a4[30][29] ),
    .B2(_03661_),
    .Y(_03850_));
 sky130_fd_sc_hd__o22a_4 _18574_ (.A1(_02577_),
    .A2(_03663_),
    .B1(_02563_),
    .B2(_03664_),
    .X(_03851_));
 sky130_fd_sc_hd__o22a_4 _18575_ (.A1(_02575_),
    .A2(_03666_),
    .B1(_02578_),
    .B2(_03667_),
    .X(_03852_));
 sky130_fd_sc_hd__and4_4 _18576_ (.A(_03849_),
    .B(_03850_),
    .C(_03851_),
    .D(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__inv_2 _18577_ (.A(\CPU_Xreg_value_a4[26][29] ),
    .Y(_03854_));
 sky130_fd_sc_hd__o22a_4 _18578_ (.A1(_03854_),
    .A2(_03671_),
    .B1(_02564_),
    .B2(_03672_),
    .X(_03855_));
 sky130_fd_sc_hd__o22a_4 _18579_ (.A1(_02580_),
    .A2(_03674_),
    .B1(_02569_),
    .B2(_03675_),
    .X(_03856_));
 sky130_fd_sc_hd__a22oi_4 _18580_ (.A1(\CPU_Xreg_value_a4[23][29] ),
    .A2(_03677_),
    .B1(\CPU_Xreg_value_a4[31][29] ),
    .B2(_03678_),
    .Y(_03857_));
 sky130_fd_sc_hd__inv_2 _18581_ (.A(\CPU_Xreg_value_a4[19][29] ),
    .Y(_03858_));
 sky130_fd_sc_hd__o22a_4 _18582_ (.A1(_03858_),
    .A2(_03681_),
    .B1(_02584_),
    .B2(_03682_),
    .X(_03859_));
 sky130_fd_sc_hd__and4_4 _18583_ (.A(_03855_),
    .B(_03856_),
    .C(_03857_),
    .D(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__o22a_4 _18584_ (.A1(_02561_),
    .A2(_03685_),
    .B1(_02583_),
    .B2(_03686_),
    .X(_03861_));
 sky130_fd_sc_hd__inv_2 _18585_ (.A(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__inv_2 _18586_ (.A(\CPU_Xreg_value_a4[25][29] ),
    .Y(_03863_));
 sky130_fd_sc_hd__a2bb2o_4 _18587_ (.A1_N(_03863_),
    .A2_N(_03690_),
    .B1(\CPU_Xreg_value_a4[24][29] ),
    .B2(_03691_),
    .X(_03864_));
 sky130_fd_sc_hd__inv_2 _18588_ (.A(\CPU_Xreg_value_a4[17][29] ),
    .Y(_03865_));
 sky130_fd_sc_hd__a2bb2o_4 _18589_ (.A1_N(_03865_),
    .A2_N(_03695_),
    .B1(\CPU_Xreg_value_a4[22][29] ),
    .B2(_03696_),
    .X(_03866_));
 sky130_fd_sc_hd__a211o_4 _18590_ (.A1(\CPU_Xreg_value_a4[13][29] ),
    .A2(_03693_),
    .B1(_02928_),
    .C1(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__inv_2 _18591_ (.A(\CPU_Xreg_value_a4[18][29] ),
    .Y(_03868_));
 sky130_fd_sc_hd__a2bb2o_4 _18592_ (.A1_N(_03868_),
    .A2_N(_03700_),
    .B1(\CPU_Xreg_value_a4[28][29] ),
    .B2(_03701_),
    .X(_03869_));
 sky130_fd_sc_hd__o22a_4 _18593_ (.A1(_02567_),
    .A2(_03703_),
    .B1(_02574_),
    .B2(_03704_),
    .X(_03870_));
 sky130_fd_sc_hd__inv_2 _18594_ (.A(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__inv_2 _18595_ (.A(\CPU_Xreg_value_a4[21][29] ),
    .Y(_03872_));
 sky130_fd_sc_hd__a2bb2o_4 _18596_ (.A1_N(_03872_),
    .A2_N(_03708_),
    .B1(\CPU_Xreg_value_a4[20][29] ),
    .B2(_03709_),
    .X(_03873_));
 sky130_fd_sc_hd__inv_2 _18597_ (.A(\CPU_Xreg_value_a4[27][29] ),
    .Y(_03874_));
 sky130_fd_sc_hd__a2bb2o_4 _18598_ (.A1_N(_03874_),
    .A2_N(_03712_),
    .B1(\CPU_Xreg_value_a4[29][29] ),
    .B2(_03713_),
    .X(_03875_));
 sky130_fd_sc_hd__or4_4 _18599_ (.A(_03869_),
    .B(_03871_),
    .C(_03873_),
    .D(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__or4_4 _18600_ (.A(_03862_),
    .B(_03864_),
    .C(_03867_),
    .D(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__inv_2 _18601_ (.A(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a32o_4 _18602_ (.A1(_03853_),
    .A2(_03860_),
    .A3(_03878_),
    .B1(_06107_),
    .B2(_03718_),
    .X(_03879_));
 sky130_fd_sc_hd__inv_2 _18603_ (.A(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__o22a_4 _18604_ (.A1(_06529_),
    .A2(_03655_),
    .B1(_03656_),
    .B2(_03880_),
    .X(\CPU_src2_value_a2[29] ));
 sky130_fd_sc_hd__o22a_4 _18605_ (.A1(_02598_),
    .A2(_02681_),
    .B1(_02609_),
    .B2(_02686_),
    .X(_03881_));
 sky130_fd_sc_hd__a22oi_4 _18606_ (.A1(\CPU_Xreg_value_a4[16][30] ),
    .A2(_02693_),
    .B1(\CPU_Xreg_value_a4[30][30] ),
    .B2(_02699_),
    .Y(_03882_));
 sky130_fd_sc_hd__o22a_4 _18607_ (.A1(_02605_),
    .A2(_02704_),
    .B1(_02591_),
    .B2(_02708_),
    .X(_03883_));
 sky130_fd_sc_hd__o22a_4 _18608_ (.A1(_02603_),
    .A2(_02712_),
    .B1(_02606_),
    .B2(_02715_),
    .X(_03884_));
 sky130_fd_sc_hd__and4_4 _18609_ (.A(_03881_),
    .B(_03882_),
    .C(_03883_),
    .D(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__inv_2 _18610_ (.A(\CPU_Xreg_value_a4[26][30] ),
    .Y(_03886_));
 sky130_fd_sc_hd__o22a_4 _18611_ (.A1(_03886_),
    .A2(_02721_),
    .B1(_02592_),
    .B2(_02724_),
    .X(_03887_));
 sky130_fd_sc_hd__o22a_4 _18612_ (.A1(_02608_),
    .A2(_02728_),
    .B1(_02597_),
    .B2(_02731_),
    .X(_03888_));
 sky130_fd_sc_hd__a22oi_4 _18613_ (.A1(\CPU_Xreg_value_a4[23][30] ),
    .A2(_02736_),
    .B1(\CPU_Xreg_value_a4[31][30] ),
    .B2(_02740_),
    .Y(_03889_));
 sky130_fd_sc_hd__inv_2 _18614_ (.A(\CPU_Xreg_value_a4[19][30] ),
    .Y(_03890_));
 sky130_fd_sc_hd__o22a_4 _18615_ (.A1(_03890_),
    .A2(_02744_),
    .B1(_02612_),
    .B2(_02747_),
    .X(_03891_));
 sky130_fd_sc_hd__and4_4 _18616_ (.A(_03887_),
    .B(_03888_),
    .C(_03889_),
    .D(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__o22a_4 _18617_ (.A1(_02589_),
    .A2(_02752_),
    .B1(_02611_),
    .B2(_02756_),
    .X(_03893_));
 sky130_fd_sc_hd__inv_2 _18618_ (.A(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__inv_2 _18619_ (.A(\CPU_Xreg_value_a4[25][30] ),
    .Y(_03895_));
 sky130_fd_sc_hd__a2bb2o_4 _18620_ (.A1_N(_03895_),
    .A2_N(_02761_),
    .B1(\CPU_Xreg_value_a4[24][30] ),
    .B2(_02765_),
    .X(_03896_));
 sky130_fd_sc_hd__inv_2 _18621_ (.A(\CPU_Xreg_value_a4[17][30] ),
    .Y(_03897_));
 sky130_fd_sc_hd__a2bb2o_4 _18622_ (.A1_N(_03897_),
    .A2_N(_02778_),
    .B1(\CPU_Xreg_value_a4[22][30] ),
    .B2(_02783_),
    .X(_03898_));
 sky130_fd_sc_hd__a211o_4 _18623_ (.A1(\CPU_Xreg_value_a4[13][30] ),
    .A2(_02771_),
    .B1(_02928_),
    .C1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__inv_2 _18624_ (.A(\CPU_Xreg_value_a4[18][30] ),
    .Y(_03900_));
 sky130_fd_sc_hd__a2bb2o_4 _18625_ (.A1_N(_03900_),
    .A2_N(_02789_),
    .B1(\CPU_Xreg_value_a4[28][30] ),
    .B2(_02793_),
    .X(_03901_));
 sky130_fd_sc_hd__o22a_4 _18626_ (.A1(_02595_),
    .A2(_02797_),
    .B1(_02602_),
    .B2(_02800_),
    .X(_03902_));
 sky130_fd_sc_hd__inv_2 _18627_ (.A(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__inv_2 _18628_ (.A(\CPU_Xreg_value_a4[21][30] ),
    .Y(_03904_));
 sky130_fd_sc_hd__a2bb2o_4 _18629_ (.A1_N(_03904_),
    .A2_N(_02805_),
    .B1(\CPU_Xreg_value_a4[20][30] ),
    .B2(_02809_),
    .X(_03905_));
 sky130_fd_sc_hd__inv_2 _18630_ (.A(\CPU_Xreg_value_a4[27][30] ),
    .Y(_03906_));
 sky130_fd_sc_hd__a2bb2o_4 _18631_ (.A1_N(_03906_),
    .A2_N(_02813_),
    .B1(\CPU_Xreg_value_a4[29][30] ),
    .B2(_02817_),
    .X(_03907_));
 sky130_fd_sc_hd__or4_4 _18632_ (.A(_03901_),
    .B(_03903_),
    .C(_03905_),
    .D(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__or4_4 _18633_ (.A(_03894_),
    .B(_03896_),
    .C(_03899_),
    .D(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__inv_2 _18634_ (.A(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__a32o_4 _18635_ (.A1(_03885_),
    .A2(_03892_),
    .A3(_03910_),
    .B1(_06106_),
    .B2(_02823_),
    .X(_03911_));
 sky130_fd_sc_hd__inv_2 _18636_ (.A(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__o22a_4 _18637_ (.A1(_06513_),
    .A2(_02669_),
    .B1(_02672_),
    .B2(_03912_),
    .X(\CPU_src2_value_a2[30] ));
 sky130_fd_sc_hd__o22a_4 _18638_ (.A1(_02626_),
    .A2(_02681_),
    .B1(_02637_),
    .B2(_02686_),
    .X(_03913_));
 sky130_fd_sc_hd__a22oi_4 _18639_ (.A1(\CPU_Xreg_value_a4[16][31] ),
    .A2(_02693_),
    .B1(\CPU_Xreg_value_a4[30][31] ),
    .B2(_02699_),
    .Y(_03914_));
 sky130_fd_sc_hd__o22a_4 _18640_ (.A1(_02633_),
    .A2(_02704_),
    .B1(_02619_),
    .B2(_02708_),
    .X(_03915_));
 sky130_fd_sc_hd__o22a_4 _18641_ (.A1(_02631_),
    .A2(_02712_),
    .B1(_02634_),
    .B2(_02715_),
    .X(_03916_));
 sky130_fd_sc_hd__and4_4 _18642_ (.A(_03913_),
    .B(_03914_),
    .C(_03915_),
    .D(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__inv_2 _18643_ (.A(\CPU_Xreg_value_a4[26][31] ),
    .Y(_03918_));
 sky130_fd_sc_hd__o22a_4 _18644_ (.A1(_03918_),
    .A2(_02721_),
    .B1(_02620_),
    .B2(_02724_),
    .X(_03919_));
 sky130_fd_sc_hd__o22a_4 _18645_ (.A1(_02636_),
    .A2(_02728_),
    .B1(_02625_),
    .B2(_02731_),
    .X(_03920_));
 sky130_fd_sc_hd__a22oi_4 _18646_ (.A1(\CPU_Xreg_value_a4[23][31] ),
    .A2(_02736_),
    .B1(\CPU_Xreg_value_a4[31][31] ),
    .B2(_02740_),
    .Y(_03921_));
 sky130_fd_sc_hd__inv_2 _18647_ (.A(\CPU_Xreg_value_a4[19][31] ),
    .Y(_03922_));
 sky130_fd_sc_hd__o22a_4 _18648_ (.A1(_03922_),
    .A2(_02744_),
    .B1(_02640_),
    .B2(_02747_),
    .X(_03923_));
 sky130_fd_sc_hd__and4_4 _18649_ (.A(_03919_),
    .B(_03920_),
    .C(_03921_),
    .D(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__o22a_4 _18650_ (.A1(_02617_),
    .A2(_02752_),
    .B1(_02639_),
    .B2(_02756_),
    .X(_03925_));
 sky130_fd_sc_hd__inv_2 _18651_ (.A(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__inv_2 _18652_ (.A(\CPU_Xreg_value_a4[25][31] ),
    .Y(_03927_));
 sky130_fd_sc_hd__a2bb2o_4 _18653_ (.A1_N(_03927_),
    .A2_N(_02761_),
    .B1(\CPU_Xreg_value_a4[24][31] ),
    .B2(_02765_),
    .X(_03928_));
 sky130_fd_sc_hd__inv_2 _18654_ (.A(\CPU_Xreg_value_a4[17][31] ),
    .Y(_03929_));
 sky130_fd_sc_hd__a2bb2o_4 _18655_ (.A1_N(_03929_),
    .A2_N(_02778_),
    .B1(\CPU_Xreg_value_a4[22][31] ),
    .B2(_02783_),
    .X(_03930_));
 sky130_fd_sc_hd__a211o_4 _18656_ (.A1(\CPU_Xreg_value_a4[13][31] ),
    .A2(_02771_),
    .B1(_02928_),
    .C1(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__inv_2 _18657_ (.A(\CPU_Xreg_value_a4[18][31] ),
    .Y(_03932_));
 sky130_fd_sc_hd__a2bb2o_4 _18658_ (.A1_N(_03932_),
    .A2_N(_02789_),
    .B1(\CPU_Xreg_value_a4[28][31] ),
    .B2(_02793_),
    .X(_03933_));
 sky130_fd_sc_hd__o22a_4 _18659_ (.A1(_02623_),
    .A2(_02797_),
    .B1(_02630_),
    .B2(_02800_),
    .X(_03934_));
 sky130_fd_sc_hd__inv_2 _18660_ (.A(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__inv_2 _18661_ (.A(\CPU_Xreg_value_a4[21][31] ),
    .Y(_03936_));
 sky130_fd_sc_hd__a2bb2o_4 _18662_ (.A1_N(_03936_),
    .A2_N(_02805_),
    .B1(\CPU_Xreg_value_a4[20][31] ),
    .B2(_02809_),
    .X(_03937_));
 sky130_fd_sc_hd__inv_2 _18663_ (.A(\CPU_Xreg_value_a4[27][31] ),
    .Y(_03938_));
 sky130_fd_sc_hd__a2bb2o_4 _18664_ (.A1_N(_03938_),
    .A2_N(_02813_),
    .B1(\CPU_Xreg_value_a4[29][31] ),
    .B2(_02817_),
    .X(_03939_));
 sky130_fd_sc_hd__or4_4 _18665_ (.A(_03933_),
    .B(_03935_),
    .C(_03937_),
    .D(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__or4_4 _18666_ (.A(_03926_),
    .B(_03928_),
    .C(_03931_),
    .D(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__inv_2 _18667_ (.A(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__a32o_4 _18668_ (.A1(_03917_),
    .A2(_03924_),
    .A3(_03942_),
    .B1(_06105_),
    .B2(_02823_),
    .X(_03943_));
 sky130_fd_sc_hd__inv_2 _18669_ (.A(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__o22a_4 _18670_ (.A1(_06501_),
    .A2(_02669_),
    .B1(_02672_),
    .B2(_03944_),
    .X(\CPU_src2_value_a2[31] ));
 sky130_fd_sc_hd__buf_2 _18671_ (.A(_04655_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_2 _18672_ (.A(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__buf_2 _18673_ (.A(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__buf_2 _18674_ (.A(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__buf_2 _18675_ (.A(_05521_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_2 _18676_ (.A(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__inv_2 _18677_ (.A(_05352_),
    .Y(_03951_));
 sky130_fd_sc_hd__buf_2 _18678_ (.A(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__buf_2 _18679_ (.A(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__a2bb2o_4 _18680_ (.A1_N(_05603_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][0] ),
    .B2(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__inv_2 _18681_ (.A(\CPU_Dmem_value_a5[8][0] ),
    .Y(_03955_));
 sky130_fd_sc_hd__buf_2 _18682_ (.A(_05434_),
    .X(_03956_));
 sky130_fd_sc_hd__buf_2 _18683_ (.A(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__inv_2 _18684_ (.A(_05856_),
    .Y(_03958_));
 sky130_fd_sc_hd__buf_2 _18685_ (.A(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__buf_2 _18686_ (.A(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__a2bb2o_4 _18687_ (.A1_N(_03955_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][0] ),
    .B2(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__inv_2 _18688_ (.A(\CPU_Dmem_value_a5[2][0] ),
    .Y(_03962_));
 sky130_fd_sc_hd__buf_2 _18689_ (.A(_04895_),
    .X(_03963_));
 sky130_fd_sc_hd__buf_2 _18690_ (.A(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__o21ai_4 _18691_ (.A1(_03962_),
    .A2(_03964_),
    .B1(_03946_),
    .Y(_03965_));
 sky130_fd_sc_hd__buf_2 _18692_ (.A(_04982_),
    .X(_03966_));
 sky130_fd_sc_hd__buf_2 _18693_ (.A(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__inv_2 _18694_ (.A(_05606_),
    .Y(_03968_));
 sky130_fd_sc_hd__buf_2 _18695_ (.A(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__buf_2 _18696_ (.A(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__a2bb2o_4 _18697_ (.A1_N(_05064_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][0] ),
    .B2(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__or4_4 _18698_ (.A(_03954_),
    .B(_03961_),
    .C(_03965_),
    .D(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__buf_2 _18699_ (.A(_04806_),
    .X(_03973_));
 sky130_fd_sc_hd__o22a_4 _18700_ (.A1(_04890_),
    .A2(_03973_),
    .B1(_05151_),
    .B2(_05068_),
    .X(_03974_));
 sky130_fd_sc_hd__buf_2 _18701_ (.A(_05239_),
    .X(_03975_));
 sky130_fd_sc_hd__inv_2 _18702_ (.A(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__inv_2 _18703_ (.A(_05689_),
    .Y(_03977_));
 sky130_fd_sc_hd__buf_2 _18704_ (.A(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__a22oi_4 _18705_ (.A1(\CPU_Dmem_value_a5[6][0] ),
    .A2(_03976_),
    .B1(\CPU_Dmem_value_a5[11][0] ),
    .B2(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__buf_2 _18706_ (.A(_05938_),
    .X(_03980_));
 sky130_fd_sc_hd__inv_2 _18707_ (.A(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__inv_2 _18708_ (.A(_05154_),
    .Y(_03982_));
 sky130_fd_sc_hd__buf_2 _18709_ (.A(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__a22oi_4 _18710_ (.A1(\CPU_Dmem_value_a5[14][0] ),
    .A2(_03981_),
    .B1(\CPU_Dmem_value_a5[5][0] ),
    .B2(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__buf_2 _18711_ (.A(_05772_),
    .X(_03985_));
 sky130_fd_sc_hd__inv_2 _18712_ (.A(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__inv_2 _18713_ (.A(_06022_),
    .Y(_03987_));
 sky130_fd_sc_hd__buf_2 _18714_ (.A(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__a22oi_4 _18715_ (.A1(\CPU_Dmem_value_a5[12][0] ),
    .A2(_03986_),
    .B1(\CPU_Dmem_value_a5[15][0] ),
    .B2(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__and4_4 _18716_ (.A(_03974_),
    .B(_03979_),
    .C(_03984_),
    .D(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__inv_2 _18717_ (.A(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__o22a_4 _18718_ (.A1(\CPU_Dmem_value_a5[0][0] ),
    .A2(_03948_),
    .B1(_03972_),
    .B2(_03991_),
    .X(\CPU_dmem_rd_data_a4[0] ));
 sky130_fd_sc_hd__inv_2 _18719_ (.A(\CPU_Dmem_value_a5[9][1] ),
    .Y(_03992_));
 sky130_fd_sc_hd__a2bb2o_4 _18720_ (.A1_N(_03992_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][1] ),
    .B2(_03953_),
    .X(_03993_));
 sky130_fd_sc_hd__inv_2 _18721_ (.A(\CPU_Dmem_value_a5[8][1] ),
    .Y(_03994_));
 sky130_fd_sc_hd__a2bb2o_4 _18722_ (.A1_N(_03994_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][1] ),
    .B2(_03960_),
    .X(_03995_));
 sky130_fd_sc_hd__o21ai_4 _18723_ (.A1(_04977_),
    .A2(_03964_),
    .B1(_03946_),
    .Y(_03996_));
 sky130_fd_sc_hd__a2bb2o_4 _18724_ (.A1_N(_05062_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][1] ),
    .B2(_03970_),
    .X(_03997_));
 sky130_fd_sc_hd__or4_4 _18725_ (.A(_03993_),
    .B(_03995_),
    .C(_03996_),
    .D(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__inv_2 _18726_ (.A(\CPU_Dmem_value_a5[1][1] ),
    .Y(_03999_));
 sky130_fd_sc_hd__buf_2 _18727_ (.A(_03973_),
    .X(_04000_));
 sky130_fd_sc_hd__inv_2 _18728_ (.A(_05068_),
    .Y(_04001_));
 sky130_fd_sc_hd__buf_2 _18729_ (.A(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__a2bb2o_4 _18730_ (.A1_N(_03999_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][1] ),
    .B2(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__buf_2 _18731_ (.A(_03975_),
    .X(_04004_));
 sky130_fd_sc_hd__a2bb2o_4 _18732_ (.A1_N(_05346_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][1] ),
    .B2(_03978_),
    .X(_04005_));
 sky130_fd_sc_hd__buf_2 _18733_ (.A(_03980_),
    .X(_04006_));
 sky130_fd_sc_hd__a2bb2o_4 _18734_ (.A1_N(_06018_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][1] ),
    .B2(_03983_),
    .X(_04007_));
 sky130_fd_sc_hd__inv_2 _18735_ (.A(\CPU_Dmem_value_a5[12][1] ),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_2 _18736_ (.A(_03985_),
    .X(_04009_));
 sky130_fd_sc_hd__a2bb2o_4 _18737_ (.A1_N(_04008_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][1] ),
    .B2(_03988_),
    .X(_04010_));
 sky130_fd_sc_hd__or4_4 _18738_ (.A(_04003_),
    .B(_04005_),
    .C(_04007_),
    .D(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__o22a_4 _18739_ (.A1(\CPU_Dmem_value_a5[0][1] ),
    .A2(_03948_),
    .B1(_03998_),
    .B2(_04011_),
    .X(\CPU_dmem_rd_data_a4[1] ));
 sky130_fd_sc_hd__inv_2 _18740_ (.A(\CPU_Dmem_value_a5[9][2] ),
    .Y(_04012_));
 sky130_fd_sc_hd__a2bb2o_4 _18741_ (.A1_N(_04012_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][2] ),
    .B2(_03953_),
    .X(_04013_));
 sky130_fd_sc_hd__inv_2 _18742_ (.A(\CPU_Dmem_value_a5[8][2] ),
    .Y(_04014_));
 sky130_fd_sc_hd__a2bb2o_4 _18743_ (.A1_N(_04014_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][2] ),
    .B2(_03960_),
    .X(_04015_));
 sky130_fd_sc_hd__inv_2 _18744_ (.A(\CPU_Dmem_value_a5[2][2] ),
    .Y(_04016_));
 sky130_fd_sc_hd__o21ai_4 _18745_ (.A1(_04016_),
    .A2(_03964_),
    .B1(_03946_),
    .Y(_04017_));
 sky130_fd_sc_hd__inv_2 _18746_ (.A(\CPU_Dmem_value_a5[3][2] ),
    .Y(_04018_));
 sky130_fd_sc_hd__a2bb2o_4 _18747_ (.A1_N(_04018_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][2] ),
    .B2(_03970_),
    .X(_04019_));
 sky130_fd_sc_hd__or4_4 _18748_ (.A(_04013_),
    .B(_04015_),
    .C(_04017_),
    .D(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__inv_2 _18749_ (.A(\CPU_Dmem_value_a5[1][2] ),
    .Y(_04021_));
 sky130_fd_sc_hd__a2bb2o_4 _18750_ (.A1_N(_04021_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][2] ),
    .B2(_04002_),
    .X(_04022_));
 sky130_fd_sc_hd__a2bb2o_4 _18751_ (.A1_N(_05344_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][2] ),
    .B2(_03978_),
    .X(_04023_));
 sky130_fd_sc_hd__a2bb2o_4 _18752_ (.A1_N(_06016_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][2] ),
    .B2(_03983_),
    .X(_04024_));
 sky130_fd_sc_hd__a2bb2o_4 _18753_ (.A1_N(_05850_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][2] ),
    .B2(_03988_),
    .X(_04025_));
 sky130_fd_sc_hd__or4_4 _18754_ (.A(_04022_),
    .B(_04023_),
    .C(_04024_),
    .D(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__o22a_4 _18755_ (.A1(\CPU_Dmem_value_a5[0][2] ),
    .A2(_03948_),
    .B1(_04020_),
    .B2(_04026_),
    .X(\CPU_dmem_rd_data_a4[2] ));
 sky130_fd_sc_hd__a2bb2o_4 _18756_ (.A1_N(_05597_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][3] ),
    .B2(_03953_),
    .X(_04027_));
 sky130_fd_sc_hd__a2bb2o_4 _18757_ (.A1_N(_05512_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][3] ),
    .B2(_03960_),
    .X(_04028_));
 sky130_fd_sc_hd__inv_2 _18758_ (.A(\CPU_Dmem_value_a5[2][3] ),
    .Y(_04029_));
 sky130_fd_sc_hd__o21ai_4 _18759_ (.A1(_04029_),
    .A2(_03964_),
    .B1(_03946_),
    .Y(_04030_));
 sky130_fd_sc_hd__inv_2 _18760_ (.A(\CPU_Dmem_value_a5[3][3] ),
    .Y(_04031_));
 sky130_fd_sc_hd__a2bb2o_4 _18761_ (.A1_N(_04031_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][3] ),
    .B2(_03970_),
    .X(_04032_));
 sky130_fd_sc_hd__or4_4 _18762_ (.A(_04027_),
    .B(_04028_),
    .C(_04030_),
    .D(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__inv_2 _18763_ (.A(\CPU_Dmem_value_a5[1][3] ),
    .Y(_04034_));
 sky130_fd_sc_hd__a2bb2o_4 _18764_ (.A1_N(_04034_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][3] ),
    .B2(_04002_),
    .X(_04035_));
 sky130_fd_sc_hd__inv_2 _18765_ (.A(\CPU_Dmem_value_a5[6][3] ),
    .Y(_04036_));
 sky130_fd_sc_hd__a2bb2o_4 _18766_ (.A1_N(_04036_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][3] ),
    .B2(_03978_),
    .X(_04037_));
 sky130_fd_sc_hd__a2bb2o_4 _18767_ (.A1_N(_06014_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][3] ),
    .B2(_03983_),
    .X(_04038_));
 sky130_fd_sc_hd__a2bb2o_4 _18768_ (.A1_N(_05848_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][3] ),
    .B2(_03988_),
    .X(_04039_));
 sky130_fd_sc_hd__or4_4 _18769_ (.A(_04035_),
    .B(_04037_),
    .C(_04038_),
    .D(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__o22a_4 _18770_ (.A1(\CPU_Dmem_value_a5[0][3] ),
    .A2(_03948_),
    .B1(_04033_),
    .B2(_04040_),
    .X(\CPU_dmem_rd_data_a4[3] ));
 sky130_fd_sc_hd__inv_2 _18771_ (.A(\CPU_Dmem_value_a5[9][4] ),
    .Y(_04041_));
 sky130_fd_sc_hd__a2bb2o_4 _18772_ (.A1_N(_04041_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][4] ),
    .B2(_03953_),
    .X(_04042_));
 sky130_fd_sc_hd__inv_2 _18773_ (.A(\CPU_Dmem_value_a5[8][4] ),
    .Y(_04043_));
 sky130_fd_sc_hd__a2bb2o_4 _18774_ (.A1_N(_04043_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][4] ),
    .B2(_03960_),
    .X(_04044_));
 sky130_fd_sc_hd__inv_2 _18775_ (.A(\CPU_Dmem_value_a5[2][4] ),
    .Y(_04045_));
 sky130_fd_sc_hd__buf_2 _18776_ (.A(_03945_),
    .X(_04046_));
 sky130_fd_sc_hd__o21ai_4 _18777_ (.A1(_04045_),
    .A2(_03964_),
    .B1(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__inv_2 _18778_ (.A(\CPU_Dmem_value_a5[3][4] ),
    .Y(_04048_));
 sky130_fd_sc_hd__a2bb2o_4 _18779_ (.A1_N(_04048_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][4] ),
    .B2(_03970_),
    .X(_04049_));
 sky130_fd_sc_hd__or4_4 _18780_ (.A(_04042_),
    .B(_04044_),
    .C(_04047_),
    .D(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__inv_2 _18781_ (.A(\CPU_Dmem_value_a5[1][4] ),
    .Y(_04051_));
 sky130_fd_sc_hd__a2bb2o_4 _18782_ (.A1_N(_04051_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][4] ),
    .B2(_04002_),
    .X(_04052_));
 sky130_fd_sc_hd__inv_2 _18783_ (.A(\CPU_Dmem_value_a5[6][4] ),
    .Y(_04053_));
 sky130_fd_sc_hd__a2bb2o_4 _18784_ (.A1_N(_04053_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][4] ),
    .B2(_03978_),
    .X(_04054_));
 sky130_fd_sc_hd__inv_2 _18785_ (.A(\CPU_Dmem_value_a5[14][4] ),
    .Y(_04055_));
 sky130_fd_sc_hd__a2bb2o_4 _18786_ (.A1_N(_04055_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][4] ),
    .B2(_03983_),
    .X(_04056_));
 sky130_fd_sc_hd__inv_2 _18787_ (.A(\CPU_Dmem_value_a5[12][4] ),
    .Y(_04057_));
 sky130_fd_sc_hd__a2bb2o_4 _18788_ (.A1_N(_04057_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][4] ),
    .B2(_03988_),
    .X(_04058_));
 sky130_fd_sc_hd__or4_4 _18789_ (.A(_04052_),
    .B(_04054_),
    .C(_04056_),
    .D(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__o22a_4 _18790_ (.A1(\CPU_Dmem_value_a5[0][4] ),
    .A2(_03948_),
    .B1(_04050_),
    .B2(_04059_),
    .X(\CPU_dmem_rd_data_a4[4] ));
 sky130_fd_sc_hd__inv_2 _18791_ (.A(\CPU_Dmem_value_a5[9][5] ),
    .Y(_04060_));
 sky130_fd_sc_hd__a2bb2o_4 _18792_ (.A1_N(_04060_),
    .A2_N(_03950_),
    .B1(\CPU_Dmem_value_a5[7][5] ),
    .B2(_03953_),
    .X(_04061_));
 sky130_fd_sc_hd__inv_2 _18793_ (.A(\CPU_Dmem_value_a5[8][5] ),
    .Y(_04062_));
 sky130_fd_sc_hd__a2bb2o_4 _18794_ (.A1_N(_04062_),
    .A2_N(_03957_),
    .B1(\CPU_Dmem_value_a5[13][5] ),
    .B2(_03960_),
    .X(_04063_));
 sky130_fd_sc_hd__inv_2 _18795_ (.A(\CPU_Dmem_value_a5[2][5] ),
    .Y(_04064_));
 sky130_fd_sc_hd__o21ai_4 _18796_ (.A1(_04064_),
    .A2(_03964_),
    .B1(_04046_),
    .Y(_04065_));
 sky130_fd_sc_hd__inv_2 _18797_ (.A(\CPU_Dmem_value_a5[3][5] ),
    .Y(_04066_));
 sky130_fd_sc_hd__a2bb2o_4 _18798_ (.A1_N(_04066_),
    .A2_N(_03967_),
    .B1(\CPU_Dmem_value_a5[10][5] ),
    .B2(_03970_),
    .X(_04067_));
 sky130_fd_sc_hd__or4_4 _18799_ (.A(_04061_),
    .B(_04063_),
    .C(_04065_),
    .D(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__inv_2 _18800_ (.A(\CPU_Dmem_value_a5[1][5] ),
    .Y(_04069_));
 sky130_fd_sc_hd__a2bb2o_4 _18801_ (.A1_N(_04069_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][5] ),
    .B2(_04002_),
    .X(_04070_));
 sky130_fd_sc_hd__inv_2 _18802_ (.A(\CPU_Dmem_value_a5[6][5] ),
    .Y(_04071_));
 sky130_fd_sc_hd__a2bb2o_4 _18803_ (.A1_N(_04071_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][5] ),
    .B2(_03978_),
    .X(_04072_));
 sky130_fd_sc_hd__inv_2 _18804_ (.A(\CPU_Dmem_value_a5[14][5] ),
    .Y(_04073_));
 sky130_fd_sc_hd__a2bb2o_4 _18805_ (.A1_N(_04073_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][5] ),
    .B2(_03983_),
    .X(_04074_));
 sky130_fd_sc_hd__inv_2 _18806_ (.A(\CPU_Dmem_value_a5[12][5] ),
    .Y(_04075_));
 sky130_fd_sc_hd__a2bb2o_4 _18807_ (.A1_N(_04075_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][5] ),
    .B2(_03988_),
    .X(_04076_));
 sky130_fd_sc_hd__or4_4 _18808_ (.A(_04070_),
    .B(_04072_),
    .C(_04074_),
    .D(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__o22a_4 _18809_ (.A1(\CPU_Dmem_value_a5[0][5] ),
    .A2(_03948_),
    .B1(_04068_),
    .B2(_04077_),
    .X(\CPU_dmem_rd_data_a4[5] ));
 sky130_fd_sc_hd__buf_2 _18810_ (.A(_03947_),
    .X(_04078_));
 sky130_fd_sc_hd__inv_2 _18811_ (.A(\CPU_Dmem_value_a5[9][6] ),
    .Y(_04079_));
 sky130_fd_sc_hd__buf_2 _18812_ (.A(_03949_),
    .X(_04080_));
 sky130_fd_sc_hd__buf_2 _18813_ (.A(_03952_),
    .X(_04081_));
 sky130_fd_sc_hd__a2bb2o_4 _18814_ (.A1_N(_04079_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][6] ),
    .B2(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__inv_2 _18815_ (.A(\CPU_Dmem_value_a5[8][6] ),
    .Y(_04083_));
 sky130_fd_sc_hd__buf_2 _18816_ (.A(_03956_),
    .X(_04084_));
 sky130_fd_sc_hd__buf_2 _18817_ (.A(_03959_),
    .X(_04085_));
 sky130_fd_sc_hd__a2bb2o_4 _18818_ (.A1_N(_04083_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][6] ),
    .B2(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__inv_2 _18819_ (.A(\CPU_Dmem_value_a5[2][6] ),
    .Y(_04087_));
 sky130_fd_sc_hd__buf_2 _18820_ (.A(_03963_),
    .X(_04088_));
 sky130_fd_sc_hd__o21ai_4 _18821_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04046_),
    .Y(_04089_));
 sky130_fd_sc_hd__inv_2 _18822_ (.A(\CPU_Dmem_value_a5[3][6] ),
    .Y(_04090_));
 sky130_fd_sc_hd__buf_2 _18823_ (.A(_03966_),
    .X(_04091_));
 sky130_fd_sc_hd__buf_2 _18824_ (.A(_03969_),
    .X(_04092_));
 sky130_fd_sc_hd__a2bb2o_4 _18825_ (.A1_N(_04090_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][6] ),
    .B2(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__or4_4 _18826_ (.A(_04082_),
    .B(_04086_),
    .C(_04089_),
    .D(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__inv_2 _18827_ (.A(\CPU_Dmem_value_a5[1][6] ),
    .Y(_04095_));
 sky130_fd_sc_hd__a2bb2o_4 _18828_ (.A1_N(_04095_),
    .A2_N(_04000_),
    .B1(\CPU_Dmem_value_a5[4][6] ),
    .B2(_04002_),
    .X(_04096_));
 sky130_fd_sc_hd__inv_2 _18829_ (.A(\CPU_Dmem_value_a5[6][6] ),
    .Y(_04097_));
 sky130_fd_sc_hd__buf_2 _18830_ (.A(_03977_),
    .X(_04098_));
 sky130_fd_sc_hd__buf_2 _18831_ (.A(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__a2bb2o_4 _18832_ (.A1_N(_04097_),
    .A2_N(_04004_),
    .B1(\CPU_Dmem_value_a5[11][6] ),
    .B2(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__inv_2 _18833_ (.A(\CPU_Dmem_value_a5[14][6] ),
    .Y(_04101_));
 sky130_fd_sc_hd__buf_2 _18834_ (.A(_03982_),
    .X(_04102_));
 sky130_fd_sc_hd__buf_2 _18835_ (.A(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__a2bb2o_4 _18836_ (.A1_N(_04101_),
    .A2_N(_04006_),
    .B1(\CPU_Dmem_value_a5[5][6] ),
    .B2(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__inv_2 _18837_ (.A(\CPU_Dmem_value_a5[12][6] ),
    .Y(_04105_));
 sky130_fd_sc_hd__buf_2 _18838_ (.A(_03987_),
    .X(_04106_));
 sky130_fd_sc_hd__buf_2 _18839_ (.A(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__a2bb2o_4 _18840_ (.A1_N(_04105_),
    .A2_N(_04009_),
    .B1(\CPU_Dmem_value_a5[15][6] ),
    .B2(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__or4_4 _18841_ (.A(_04096_),
    .B(_04100_),
    .C(_04104_),
    .D(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__o22a_4 _18842_ (.A1(\CPU_Dmem_value_a5[0][6] ),
    .A2(_04078_),
    .B1(_04094_),
    .B2(_04109_),
    .X(\CPU_dmem_rd_data_a4[6] ));
 sky130_fd_sc_hd__inv_2 _18843_ (.A(\CPU_Dmem_value_a5[9][7] ),
    .Y(_04110_));
 sky130_fd_sc_hd__a2bb2o_4 _18844_ (.A1_N(_04110_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][7] ),
    .B2(_04081_),
    .X(_04111_));
 sky130_fd_sc_hd__inv_2 _18845_ (.A(\CPU_Dmem_value_a5[8][7] ),
    .Y(_04112_));
 sky130_fd_sc_hd__a2bb2o_4 _18846_ (.A1_N(_04112_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][7] ),
    .B2(_04085_),
    .X(_04113_));
 sky130_fd_sc_hd__inv_2 _18847_ (.A(\CPU_Dmem_value_a5[2][7] ),
    .Y(_04114_));
 sky130_fd_sc_hd__o21ai_4 _18848_ (.A1(_04114_),
    .A2(_04088_),
    .B1(_04046_),
    .Y(_04115_));
 sky130_fd_sc_hd__inv_2 _18849_ (.A(\CPU_Dmem_value_a5[3][7] ),
    .Y(_04116_));
 sky130_fd_sc_hd__a2bb2o_4 _18850_ (.A1_N(_04116_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][7] ),
    .B2(_04092_),
    .X(_04117_));
 sky130_fd_sc_hd__or4_4 _18851_ (.A(_04111_),
    .B(_04113_),
    .C(_04115_),
    .D(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__inv_2 _18852_ (.A(\CPU_Dmem_value_a5[1][7] ),
    .Y(_04119_));
 sky130_fd_sc_hd__buf_2 _18853_ (.A(_03973_),
    .X(_04120_));
 sky130_fd_sc_hd__buf_2 _18854_ (.A(_04001_),
    .X(_04121_));
 sky130_fd_sc_hd__a2bb2o_4 _18855_ (.A1_N(_04119_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][7] ),
    .B2(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__inv_2 _18856_ (.A(\CPU_Dmem_value_a5[6][7] ),
    .Y(_04123_));
 sky130_fd_sc_hd__buf_2 _18857_ (.A(_03975_),
    .X(_04124_));
 sky130_fd_sc_hd__a2bb2o_4 _18858_ (.A1_N(_04123_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][7] ),
    .B2(_04099_),
    .X(_04125_));
 sky130_fd_sc_hd__inv_2 _18859_ (.A(\CPU_Dmem_value_a5[14][7] ),
    .Y(_04126_));
 sky130_fd_sc_hd__buf_2 _18860_ (.A(_03980_),
    .X(_04127_));
 sky130_fd_sc_hd__a2bb2o_4 _18861_ (.A1_N(_04126_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][7] ),
    .B2(_04103_),
    .X(_04128_));
 sky130_fd_sc_hd__inv_2 _18862_ (.A(\CPU_Dmem_value_a5[12][7] ),
    .Y(_04129_));
 sky130_fd_sc_hd__buf_2 _18863_ (.A(_03985_),
    .X(_04130_));
 sky130_fd_sc_hd__a2bb2o_4 _18864_ (.A1_N(_04129_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][7] ),
    .B2(_04107_),
    .X(_04131_));
 sky130_fd_sc_hd__or4_4 _18865_ (.A(_04122_),
    .B(_04125_),
    .C(_04128_),
    .D(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__o22a_4 _18866_ (.A1(\CPU_Dmem_value_a5[0][7] ),
    .A2(_04078_),
    .B1(_04118_),
    .B2(_04132_),
    .X(\CPU_dmem_rd_data_a4[7] ));
 sky130_fd_sc_hd__inv_2 _18867_ (.A(\CPU_Dmem_value_a5[9][8] ),
    .Y(_04133_));
 sky130_fd_sc_hd__a2bb2o_4 _18868_ (.A1_N(_04133_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][8] ),
    .B2(_04081_),
    .X(_04134_));
 sky130_fd_sc_hd__inv_2 _18869_ (.A(\CPU_Dmem_value_a5[8][8] ),
    .Y(_04135_));
 sky130_fd_sc_hd__a2bb2o_4 _18870_ (.A1_N(_04135_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][8] ),
    .B2(_04085_),
    .X(_04136_));
 sky130_fd_sc_hd__inv_2 _18871_ (.A(\CPU_Dmem_value_a5[2][8] ),
    .Y(_04137_));
 sky130_fd_sc_hd__o21ai_4 _18872_ (.A1(_04137_),
    .A2(_04088_),
    .B1(_04046_),
    .Y(_04138_));
 sky130_fd_sc_hd__inv_2 _18873_ (.A(\CPU_Dmem_value_a5[3][8] ),
    .Y(_04139_));
 sky130_fd_sc_hd__a2bb2o_4 _18874_ (.A1_N(_04139_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][8] ),
    .B2(_04092_),
    .X(_04140_));
 sky130_fd_sc_hd__or4_4 _18875_ (.A(_04134_),
    .B(_04136_),
    .C(_04138_),
    .D(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__inv_2 _18876_ (.A(\CPU_Dmem_value_a5[1][8] ),
    .Y(_04142_));
 sky130_fd_sc_hd__a2bb2o_4 _18877_ (.A1_N(_04142_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][8] ),
    .B2(_04121_),
    .X(_04143_));
 sky130_fd_sc_hd__inv_2 _18878_ (.A(\CPU_Dmem_value_a5[6][8] ),
    .Y(_04144_));
 sky130_fd_sc_hd__a2bb2o_4 _18879_ (.A1_N(_04144_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][8] ),
    .B2(_04099_),
    .X(_04145_));
 sky130_fd_sc_hd__inv_2 _18880_ (.A(\CPU_Dmem_value_a5[14][8] ),
    .Y(_04146_));
 sky130_fd_sc_hd__a2bb2o_4 _18881_ (.A1_N(_04146_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][8] ),
    .B2(_04103_),
    .X(_04147_));
 sky130_fd_sc_hd__inv_2 _18882_ (.A(\CPU_Dmem_value_a5[12][8] ),
    .Y(_04148_));
 sky130_fd_sc_hd__a2bb2o_4 _18883_ (.A1_N(_04148_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][8] ),
    .B2(_04107_),
    .X(_04149_));
 sky130_fd_sc_hd__or4_4 _18884_ (.A(_04143_),
    .B(_04145_),
    .C(_04147_),
    .D(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__o22a_4 _18885_ (.A1(\CPU_Dmem_value_a5[0][8] ),
    .A2(_04078_),
    .B1(_04141_),
    .B2(_04150_),
    .X(\CPU_dmem_rd_data_a4[8] ));
 sky130_fd_sc_hd__inv_2 _18886_ (.A(\CPU_Dmem_value_a5[9][9] ),
    .Y(_04151_));
 sky130_fd_sc_hd__a2bb2o_4 _18887_ (.A1_N(_04151_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][9] ),
    .B2(_04081_),
    .X(_04152_));
 sky130_fd_sc_hd__inv_2 _18888_ (.A(\CPU_Dmem_value_a5[8][9] ),
    .Y(_04153_));
 sky130_fd_sc_hd__a2bb2o_4 _18889_ (.A1_N(_04153_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][9] ),
    .B2(_04085_),
    .X(_04154_));
 sky130_fd_sc_hd__inv_2 _18890_ (.A(\CPU_Dmem_value_a5[2][9] ),
    .Y(_04155_));
 sky130_fd_sc_hd__o21ai_4 _18891_ (.A1(_04155_),
    .A2(_04088_),
    .B1(_04046_),
    .Y(_04156_));
 sky130_fd_sc_hd__inv_2 _18892_ (.A(\CPU_Dmem_value_a5[3][9] ),
    .Y(_04157_));
 sky130_fd_sc_hd__a2bb2o_4 _18893_ (.A1_N(_04157_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][9] ),
    .B2(_04092_),
    .X(_04158_));
 sky130_fd_sc_hd__or4_4 _18894_ (.A(_04152_),
    .B(_04154_),
    .C(_04156_),
    .D(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__inv_2 _18895_ (.A(\CPU_Dmem_value_a5[1][9] ),
    .Y(_04160_));
 sky130_fd_sc_hd__a2bb2o_4 _18896_ (.A1_N(_04160_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][9] ),
    .B2(_04121_),
    .X(_04161_));
 sky130_fd_sc_hd__inv_2 _18897_ (.A(\CPU_Dmem_value_a5[6][9] ),
    .Y(_04162_));
 sky130_fd_sc_hd__a2bb2o_4 _18898_ (.A1_N(_04162_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][9] ),
    .B2(_04099_),
    .X(_04163_));
 sky130_fd_sc_hd__inv_2 _18899_ (.A(\CPU_Dmem_value_a5[14][9] ),
    .Y(_04164_));
 sky130_fd_sc_hd__a2bb2o_4 _18900_ (.A1_N(_04164_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][9] ),
    .B2(_04103_),
    .X(_04165_));
 sky130_fd_sc_hd__inv_2 _18901_ (.A(\CPU_Dmem_value_a5[12][9] ),
    .Y(_04166_));
 sky130_fd_sc_hd__a2bb2o_4 _18902_ (.A1_N(_04166_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][9] ),
    .B2(_04107_),
    .X(_04167_));
 sky130_fd_sc_hd__or4_4 _18903_ (.A(_04161_),
    .B(_04163_),
    .C(_04165_),
    .D(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__o22a_4 _18904_ (.A1(\CPU_Dmem_value_a5[0][9] ),
    .A2(_04078_),
    .B1(_04159_),
    .B2(_04168_),
    .X(\CPU_dmem_rd_data_a4[9] ));
 sky130_fd_sc_hd__inv_2 _18905_ (.A(\CPU_Dmem_value_a5[9][10] ),
    .Y(_04169_));
 sky130_fd_sc_hd__a2bb2o_4 _18906_ (.A1_N(_04169_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][10] ),
    .B2(_04081_),
    .X(_04170_));
 sky130_fd_sc_hd__inv_2 _18907_ (.A(\CPU_Dmem_value_a5[8][10] ),
    .Y(_04171_));
 sky130_fd_sc_hd__a2bb2o_4 _18908_ (.A1_N(_04171_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][10] ),
    .B2(_04085_),
    .X(_04172_));
 sky130_fd_sc_hd__inv_2 _18909_ (.A(\CPU_Dmem_value_a5[2][10] ),
    .Y(_04173_));
 sky130_fd_sc_hd__buf_2 _18910_ (.A(_04655_),
    .X(_04174_));
 sky130_fd_sc_hd__o21ai_4 _18911_ (.A1(_04173_),
    .A2(_04088_),
    .B1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__inv_2 _18912_ (.A(\CPU_Dmem_value_a5[3][10] ),
    .Y(_04176_));
 sky130_fd_sc_hd__a2bb2o_4 _18913_ (.A1_N(_04176_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][10] ),
    .B2(_04092_),
    .X(_04177_));
 sky130_fd_sc_hd__or4_4 _18914_ (.A(_04170_),
    .B(_04172_),
    .C(_04175_),
    .D(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__inv_2 _18915_ (.A(\CPU_Dmem_value_a5[1][10] ),
    .Y(_04179_));
 sky130_fd_sc_hd__a2bb2o_4 _18916_ (.A1_N(_04179_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][10] ),
    .B2(_04121_),
    .X(_04180_));
 sky130_fd_sc_hd__inv_2 _18917_ (.A(\CPU_Dmem_value_a5[6][10] ),
    .Y(_04181_));
 sky130_fd_sc_hd__a2bb2o_4 _18918_ (.A1_N(_04181_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][10] ),
    .B2(_04099_),
    .X(_04182_));
 sky130_fd_sc_hd__inv_2 _18919_ (.A(\CPU_Dmem_value_a5[14][10] ),
    .Y(_04183_));
 sky130_fd_sc_hd__a2bb2o_4 _18920_ (.A1_N(_04183_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][10] ),
    .B2(_04103_),
    .X(_04184_));
 sky130_fd_sc_hd__inv_2 _18921_ (.A(\CPU_Dmem_value_a5[12][10] ),
    .Y(_04185_));
 sky130_fd_sc_hd__a2bb2o_4 _18922_ (.A1_N(_04185_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][10] ),
    .B2(_04107_),
    .X(_04186_));
 sky130_fd_sc_hd__or4_4 _18923_ (.A(_04180_),
    .B(_04182_),
    .C(_04184_),
    .D(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__o22a_4 _18924_ (.A1(\CPU_Dmem_value_a5[0][10] ),
    .A2(_04078_),
    .B1(_04178_),
    .B2(_04187_),
    .X(\CPU_dmem_rd_data_a4[10] ));
 sky130_fd_sc_hd__inv_2 _18925_ (.A(\CPU_Dmem_value_a5[9][11] ),
    .Y(_04188_));
 sky130_fd_sc_hd__a2bb2o_4 _18926_ (.A1_N(_04188_),
    .A2_N(_04080_),
    .B1(\CPU_Dmem_value_a5[7][11] ),
    .B2(_04081_),
    .X(_04189_));
 sky130_fd_sc_hd__inv_2 _18927_ (.A(\CPU_Dmem_value_a5[8][11] ),
    .Y(_04190_));
 sky130_fd_sc_hd__a2bb2o_4 _18928_ (.A1_N(_04190_),
    .A2_N(_04084_),
    .B1(\CPU_Dmem_value_a5[13][11] ),
    .B2(_04085_),
    .X(_04191_));
 sky130_fd_sc_hd__inv_2 _18929_ (.A(\CPU_Dmem_value_a5[2][11] ),
    .Y(_04192_));
 sky130_fd_sc_hd__o21ai_4 _18930_ (.A1(_04192_),
    .A2(_04088_),
    .B1(_04174_),
    .Y(_04193_));
 sky130_fd_sc_hd__inv_2 _18931_ (.A(\CPU_Dmem_value_a5[3][11] ),
    .Y(_04194_));
 sky130_fd_sc_hd__a2bb2o_4 _18932_ (.A1_N(_04194_),
    .A2_N(_04091_),
    .B1(\CPU_Dmem_value_a5[10][11] ),
    .B2(_04092_),
    .X(_04195_));
 sky130_fd_sc_hd__or4_4 _18933_ (.A(_04189_),
    .B(_04191_),
    .C(_04193_),
    .D(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__inv_2 _18934_ (.A(\CPU_Dmem_value_a5[1][11] ),
    .Y(_04197_));
 sky130_fd_sc_hd__a2bb2o_4 _18935_ (.A1_N(_04197_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][11] ),
    .B2(_04121_),
    .X(_04198_));
 sky130_fd_sc_hd__inv_2 _18936_ (.A(\CPU_Dmem_value_a5[6][11] ),
    .Y(_04199_));
 sky130_fd_sc_hd__a2bb2o_4 _18937_ (.A1_N(_04199_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][11] ),
    .B2(_04099_),
    .X(_04200_));
 sky130_fd_sc_hd__inv_2 _18938_ (.A(\CPU_Dmem_value_a5[14][11] ),
    .Y(_04201_));
 sky130_fd_sc_hd__a2bb2o_4 _18939_ (.A1_N(_04201_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][11] ),
    .B2(_04103_),
    .X(_04202_));
 sky130_fd_sc_hd__inv_2 _18940_ (.A(\CPU_Dmem_value_a5[12][11] ),
    .Y(_04203_));
 sky130_fd_sc_hd__a2bb2o_4 _18941_ (.A1_N(_04203_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][11] ),
    .B2(_04107_),
    .X(_04204_));
 sky130_fd_sc_hd__or4_4 _18942_ (.A(_04198_),
    .B(_04200_),
    .C(_04202_),
    .D(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__o22a_4 _18943_ (.A1(\CPU_Dmem_value_a5[0][11] ),
    .A2(_04078_),
    .B1(_04196_),
    .B2(_04205_),
    .X(\CPU_dmem_rd_data_a4[11] ));
 sky130_fd_sc_hd__buf_2 _18944_ (.A(_03947_),
    .X(_04206_));
 sky130_fd_sc_hd__inv_2 _18945_ (.A(\CPU_Dmem_value_a5[9][12] ),
    .Y(_04207_));
 sky130_fd_sc_hd__buf_2 _18946_ (.A(_03949_),
    .X(_04208_));
 sky130_fd_sc_hd__buf_2 _18947_ (.A(_03952_),
    .X(_04209_));
 sky130_fd_sc_hd__a2bb2o_4 _18948_ (.A1_N(_04207_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][12] ),
    .B2(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__inv_2 _18949_ (.A(\CPU_Dmem_value_a5[8][12] ),
    .Y(_04211_));
 sky130_fd_sc_hd__buf_2 _18950_ (.A(_03956_),
    .X(_04212_));
 sky130_fd_sc_hd__buf_2 _18951_ (.A(_03959_),
    .X(_04213_));
 sky130_fd_sc_hd__a2bb2o_4 _18952_ (.A1_N(_04211_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][12] ),
    .B2(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__inv_2 _18953_ (.A(\CPU_Dmem_value_a5[2][12] ),
    .Y(_04215_));
 sky130_fd_sc_hd__buf_2 _18954_ (.A(_03963_),
    .X(_04216_));
 sky130_fd_sc_hd__o21ai_4 _18955_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04174_),
    .Y(_04217_));
 sky130_fd_sc_hd__inv_2 _18956_ (.A(\CPU_Dmem_value_a5[3][12] ),
    .Y(_04218_));
 sky130_fd_sc_hd__buf_2 _18957_ (.A(_03966_),
    .X(_04219_));
 sky130_fd_sc_hd__buf_2 _18958_ (.A(_03969_),
    .X(_04220_));
 sky130_fd_sc_hd__a2bb2o_4 _18959_ (.A1_N(_04218_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][12] ),
    .B2(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__or4_4 _18960_ (.A(_04210_),
    .B(_04214_),
    .C(_04217_),
    .D(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__inv_2 _18961_ (.A(\CPU_Dmem_value_a5[1][12] ),
    .Y(_04223_));
 sky130_fd_sc_hd__a2bb2o_4 _18962_ (.A1_N(_04223_),
    .A2_N(_04120_),
    .B1(\CPU_Dmem_value_a5[4][12] ),
    .B2(_04121_),
    .X(_04224_));
 sky130_fd_sc_hd__inv_2 _18963_ (.A(\CPU_Dmem_value_a5[6][12] ),
    .Y(_04225_));
 sky130_fd_sc_hd__buf_2 _18964_ (.A(_04098_),
    .X(_04226_));
 sky130_fd_sc_hd__a2bb2o_4 _18965_ (.A1_N(_04225_),
    .A2_N(_04124_),
    .B1(\CPU_Dmem_value_a5[11][12] ),
    .B2(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__inv_2 _18966_ (.A(\CPU_Dmem_value_a5[14][12] ),
    .Y(_04228_));
 sky130_fd_sc_hd__buf_2 _18967_ (.A(_04102_),
    .X(_04229_));
 sky130_fd_sc_hd__a2bb2o_4 _18968_ (.A1_N(_04228_),
    .A2_N(_04127_),
    .B1(\CPU_Dmem_value_a5[5][12] ),
    .B2(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__inv_2 _18969_ (.A(\CPU_Dmem_value_a5[12][12] ),
    .Y(_04231_));
 sky130_fd_sc_hd__buf_2 _18970_ (.A(_04106_),
    .X(_04232_));
 sky130_fd_sc_hd__a2bb2o_4 _18971_ (.A1_N(_04231_),
    .A2_N(_04130_),
    .B1(\CPU_Dmem_value_a5[15][12] ),
    .B2(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__or4_4 _18972_ (.A(_04224_),
    .B(_04227_),
    .C(_04230_),
    .D(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__o22a_4 _18973_ (.A1(\CPU_Dmem_value_a5[0][12] ),
    .A2(_04206_),
    .B1(_04222_),
    .B2(_04234_),
    .X(\CPU_dmem_rd_data_a4[12] ));
 sky130_fd_sc_hd__inv_2 _18974_ (.A(\CPU_Dmem_value_a5[9][13] ),
    .Y(_04235_));
 sky130_fd_sc_hd__a2bb2o_4 _18975_ (.A1_N(_04235_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][13] ),
    .B2(_04209_),
    .X(_04236_));
 sky130_fd_sc_hd__inv_2 _18976_ (.A(\CPU_Dmem_value_a5[8][13] ),
    .Y(_04237_));
 sky130_fd_sc_hd__a2bb2o_4 _18977_ (.A1_N(_04237_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][13] ),
    .B2(_04213_),
    .X(_04238_));
 sky130_fd_sc_hd__inv_2 _18978_ (.A(\CPU_Dmem_value_a5[2][13] ),
    .Y(_04239_));
 sky130_fd_sc_hd__o21ai_4 _18979_ (.A1(_04239_),
    .A2(_04216_),
    .B1(_04174_),
    .Y(_04240_));
 sky130_fd_sc_hd__inv_2 _18980_ (.A(\CPU_Dmem_value_a5[3][13] ),
    .Y(_04241_));
 sky130_fd_sc_hd__a2bb2o_4 _18981_ (.A1_N(_04241_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][13] ),
    .B2(_04220_),
    .X(_04242_));
 sky130_fd_sc_hd__or4_4 _18982_ (.A(_04236_),
    .B(_04238_),
    .C(_04240_),
    .D(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__inv_2 _18983_ (.A(\CPU_Dmem_value_a5[1][13] ),
    .Y(_04244_));
 sky130_fd_sc_hd__buf_2 _18984_ (.A(_03973_),
    .X(_04245_));
 sky130_fd_sc_hd__buf_2 _18985_ (.A(_04001_),
    .X(_04246_));
 sky130_fd_sc_hd__a2bb2o_4 _18986_ (.A1_N(_04244_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][13] ),
    .B2(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__inv_2 _18987_ (.A(\CPU_Dmem_value_a5[6][13] ),
    .Y(_04248_));
 sky130_fd_sc_hd__buf_2 _18988_ (.A(_03975_),
    .X(_04249_));
 sky130_fd_sc_hd__a2bb2o_4 _18989_ (.A1_N(_04248_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][13] ),
    .B2(_04226_),
    .X(_04250_));
 sky130_fd_sc_hd__inv_2 _18990_ (.A(\CPU_Dmem_value_a5[14][13] ),
    .Y(_04251_));
 sky130_fd_sc_hd__buf_2 _18991_ (.A(_03980_),
    .X(_04252_));
 sky130_fd_sc_hd__a2bb2o_4 _18992_ (.A1_N(_04251_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][13] ),
    .B2(_04229_),
    .X(_04253_));
 sky130_fd_sc_hd__inv_2 _18993_ (.A(\CPU_Dmem_value_a5[12][13] ),
    .Y(_04254_));
 sky130_fd_sc_hd__buf_2 _18994_ (.A(_03985_),
    .X(_04255_));
 sky130_fd_sc_hd__a2bb2o_4 _18995_ (.A1_N(_04254_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][13] ),
    .B2(_04232_),
    .X(_04256_));
 sky130_fd_sc_hd__or4_4 _18996_ (.A(_04247_),
    .B(_04250_),
    .C(_04253_),
    .D(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__o22a_4 _18997_ (.A1(\CPU_Dmem_value_a5[0][13] ),
    .A2(_04206_),
    .B1(_04243_),
    .B2(_04257_),
    .X(\CPU_dmem_rd_data_a4[13] ));
 sky130_fd_sc_hd__inv_2 _18998_ (.A(\CPU_Dmem_value_a5[9][14] ),
    .Y(_04258_));
 sky130_fd_sc_hd__a2bb2o_4 _18999_ (.A1_N(_04258_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][14] ),
    .B2(_04209_),
    .X(_04259_));
 sky130_fd_sc_hd__inv_2 _19000_ (.A(\CPU_Dmem_value_a5[8][14] ),
    .Y(_04260_));
 sky130_fd_sc_hd__a2bb2o_4 _19001_ (.A1_N(_04260_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][14] ),
    .B2(_04213_),
    .X(_04261_));
 sky130_fd_sc_hd__inv_2 _19002_ (.A(\CPU_Dmem_value_a5[2][14] ),
    .Y(_04262_));
 sky130_fd_sc_hd__o21ai_4 _19003_ (.A1(_04262_),
    .A2(_04216_),
    .B1(_04174_),
    .Y(_04263_));
 sky130_fd_sc_hd__inv_2 _19004_ (.A(\CPU_Dmem_value_a5[3][14] ),
    .Y(_04264_));
 sky130_fd_sc_hd__a2bb2o_4 _19005_ (.A1_N(_04264_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][14] ),
    .B2(_04220_),
    .X(_04265_));
 sky130_fd_sc_hd__or4_4 _19006_ (.A(_04259_),
    .B(_04261_),
    .C(_04263_),
    .D(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__inv_2 _19007_ (.A(\CPU_Dmem_value_a5[1][14] ),
    .Y(_04267_));
 sky130_fd_sc_hd__a2bb2o_4 _19008_ (.A1_N(_04267_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][14] ),
    .B2(_04246_),
    .X(_04268_));
 sky130_fd_sc_hd__inv_2 _19009_ (.A(\CPU_Dmem_value_a5[6][14] ),
    .Y(_04269_));
 sky130_fd_sc_hd__a2bb2o_4 _19010_ (.A1_N(_04269_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][14] ),
    .B2(_04226_),
    .X(_04270_));
 sky130_fd_sc_hd__inv_2 _19011_ (.A(\CPU_Dmem_value_a5[14][14] ),
    .Y(_04271_));
 sky130_fd_sc_hd__a2bb2o_4 _19012_ (.A1_N(_04271_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][14] ),
    .B2(_04229_),
    .X(_04272_));
 sky130_fd_sc_hd__inv_2 _19013_ (.A(\CPU_Dmem_value_a5[12][14] ),
    .Y(_04273_));
 sky130_fd_sc_hd__a2bb2o_4 _19014_ (.A1_N(_04273_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][14] ),
    .B2(_04232_),
    .X(_04274_));
 sky130_fd_sc_hd__or4_4 _19015_ (.A(_04268_),
    .B(_04270_),
    .C(_04272_),
    .D(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__o22a_4 _19016_ (.A1(\CPU_Dmem_value_a5[0][14] ),
    .A2(_04206_),
    .B1(_04266_),
    .B2(_04275_),
    .X(\CPU_dmem_rd_data_a4[14] ));
 sky130_fd_sc_hd__inv_2 _19017_ (.A(\CPU_Dmem_value_a5[9][15] ),
    .Y(_04276_));
 sky130_fd_sc_hd__a2bb2o_4 _19018_ (.A1_N(_04276_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][15] ),
    .B2(_04209_),
    .X(_04277_));
 sky130_fd_sc_hd__inv_2 _19019_ (.A(\CPU_Dmem_value_a5[8][15] ),
    .Y(_04278_));
 sky130_fd_sc_hd__a2bb2o_4 _19020_ (.A1_N(_04278_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][15] ),
    .B2(_04213_),
    .X(_04279_));
 sky130_fd_sc_hd__inv_2 _19021_ (.A(\CPU_Dmem_value_a5[2][15] ),
    .Y(_04280_));
 sky130_fd_sc_hd__o21ai_4 _19022_ (.A1(_04280_),
    .A2(_04216_),
    .B1(_04174_),
    .Y(_04281_));
 sky130_fd_sc_hd__inv_2 _19023_ (.A(\CPU_Dmem_value_a5[3][15] ),
    .Y(_04282_));
 sky130_fd_sc_hd__a2bb2o_4 _19024_ (.A1_N(_04282_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][15] ),
    .B2(_04220_),
    .X(_04283_));
 sky130_fd_sc_hd__or4_4 _19025_ (.A(_04277_),
    .B(_04279_),
    .C(_04281_),
    .D(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__inv_2 _19026_ (.A(\CPU_Dmem_value_a5[1][15] ),
    .Y(_04285_));
 sky130_fd_sc_hd__a2bb2o_4 _19027_ (.A1_N(_04285_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][15] ),
    .B2(_04246_),
    .X(_04286_));
 sky130_fd_sc_hd__inv_2 _19028_ (.A(\CPU_Dmem_value_a5[6][15] ),
    .Y(_04287_));
 sky130_fd_sc_hd__a2bb2o_4 _19029_ (.A1_N(_04287_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][15] ),
    .B2(_04226_),
    .X(_04288_));
 sky130_fd_sc_hd__inv_2 _19030_ (.A(\CPU_Dmem_value_a5[14][15] ),
    .Y(_04289_));
 sky130_fd_sc_hd__a2bb2o_4 _19031_ (.A1_N(_04289_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][15] ),
    .B2(_04229_),
    .X(_04290_));
 sky130_fd_sc_hd__inv_2 _19032_ (.A(\CPU_Dmem_value_a5[12][15] ),
    .Y(_04291_));
 sky130_fd_sc_hd__a2bb2o_4 _19033_ (.A1_N(_04291_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][15] ),
    .B2(_04232_),
    .X(_04292_));
 sky130_fd_sc_hd__or4_4 _19034_ (.A(_04286_),
    .B(_04288_),
    .C(_04290_),
    .D(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__o22a_4 _19035_ (.A1(\CPU_Dmem_value_a5[0][15] ),
    .A2(_04206_),
    .B1(_04284_),
    .B2(_04293_),
    .X(\CPU_dmem_rd_data_a4[15] ));
 sky130_fd_sc_hd__inv_2 _19036_ (.A(\CPU_Dmem_value_a5[9][16] ),
    .Y(_04294_));
 sky130_fd_sc_hd__a2bb2o_4 _19037_ (.A1_N(_04294_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][16] ),
    .B2(_04209_),
    .X(_04295_));
 sky130_fd_sc_hd__inv_2 _19038_ (.A(\CPU_Dmem_value_a5[8][16] ),
    .Y(_04296_));
 sky130_fd_sc_hd__a2bb2o_4 _19039_ (.A1_N(_04296_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][16] ),
    .B2(_04213_),
    .X(_04297_));
 sky130_fd_sc_hd__inv_2 _19040_ (.A(\CPU_Dmem_value_a5[2][16] ),
    .Y(_04298_));
 sky130_fd_sc_hd__buf_2 _19041_ (.A(_04655_),
    .X(_04299_));
 sky130_fd_sc_hd__o21ai_4 _19042_ (.A1(_04298_),
    .A2(_04216_),
    .B1(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__inv_2 _19043_ (.A(\CPU_Dmem_value_a5[3][16] ),
    .Y(_04301_));
 sky130_fd_sc_hd__a2bb2o_4 _19044_ (.A1_N(_04301_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][16] ),
    .B2(_04220_),
    .X(_04302_));
 sky130_fd_sc_hd__or4_4 _19045_ (.A(_04295_),
    .B(_04297_),
    .C(_04300_),
    .D(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__inv_2 _19046_ (.A(\CPU_Dmem_value_a5[1][16] ),
    .Y(_04304_));
 sky130_fd_sc_hd__a2bb2o_4 _19047_ (.A1_N(_04304_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][16] ),
    .B2(_04246_),
    .X(_04305_));
 sky130_fd_sc_hd__inv_2 _19048_ (.A(\CPU_Dmem_value_a5[6][16] ),
    .Y(_04306_));
 sky130_fd_sc_hd__a2bb2o_4 _19049_ (.A1_N(_04306_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][16] ),
    .B2(_04226_),
    .X(_04307_));
 sky130_fd_sc_hd__inv_2 _19050_ (.A(\CPU_Dmem_value_a5[14][16] ),
    .Y(_04308_));
 sky130_fd_sc_hd__a2bb2o_4 _19051_ (.A1_N(_04308_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][16] ),
    .B2(_04229_),
    .X(_04309_));
 sky130_fd_sc_hd__inv_2 _19052_ (.A(\CPU_Dmem_value_a5[12][16] ),
    .Y(_04310_));
 sky130_fd_sc_hd__a2bb2o_4 _19053_ (.A1_N(_04310_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][16] ),
    .B2(_04232_),
    .X(_04311_));
 sky130_fd_sc_hd__or4_4 _19054_ (.A(_04305_),
    .B(_04307_),
    .C(_04309_),
    .D(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__o22a_4 _19055_ (.A1(\CPU_Dmem_value_a5[0][16] ),
    .A2(_04206_),
    .B1(_04303_),
    .B2(_04312_),
    .X(\CPU_dmem_rd_data_a4[16] ));
 sky130_fd_sc_hd__inv_2 _19056_ (.A(\CPU_Dmem_value_a5[9][17] ),
    .Y(_04313_));
 sky130_fd_sc_hd__a2bb2o_4 _19057_ (.A1_N(_04313_),
    .A2_N(_04208_),
    .B1(\CPU_Dmem_value_a5[7][17] ),
    .B2(_04209_),
    .X(_04314_));
 sky130_fd_sc_hd__inv_2 _19058_ (.A(\CPU_Dmem_value_a5[8][17] ),
    .Y(_04315_));
 sky130_fd_sc_hd__a2bb2o_4 _19059_ (.A1_N(_04315_),
    .A2_N(_04212_),
    .B1(\CPU_Dmem_value_a5[13][17] ),
    .B2(_04213_),
    .X(_04316_));
 sky130_fd_sc_hd__inv_2 _19060_ (.A(\CPU_Dmem_value_a5[2][17] ),
    .Y(_04317_));
 sky130_fd_sc_hd__o21ai_4 _19061_ (.A1(_04317_),
    .A2(_04216_),
    .B1(_04299_),
    .Y(_04318_));
 sky130_fd_sc_hd__inv_2 _19062_ (.A(\CPU_Dmem_value_a5[3][17] ),
    .Y(_04319_));
 sky130_fd_sc_hd__a2bb2o_4 _19063_ (.A1_N(_04319_),
    .A2_N(_04219_),
    .B1(\CPU_Dmem_value_a5[10][17] ),
    .B2(_04220_),
    .X(_04320_));
 sky130_fd_sc_hd__or4_4 _19064_ (.A(_04314_),
    .B(_04316_),
    .C(_04318_),
    .D(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__inv_2 _19065_ (.A(\CPU_Dmem_value_a5[1][17] ),
    .Y(_04322_));
 sky130_fd_sc_hd__a2bb2o_4 _19066_ (.A1_N(_04322_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][17] ),
    .B2(_04246_),
    .X(_04323_));
 sky130_fd_sc_hd__inv_2 _19067_ (.A(\CPU_Dmem_value_a5[6][17] ),
    .Y(_04324_));
 sky130_fd_sc_hd__a2bb2o_4 _19068_ (.A1_N(_04324_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][17] ),
    .B2(_04226_),
    .X(_04325_));
 sky130_fd_sc_hd__inv_2 _19069_ (.A(\CPU_Dmem_value_a5[14][17] ),
    .Y(_04326_));
 sky130_fd_sc_hd__a2bb2o_4 _19070_ (.A1_N(_04326_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][17] ),
    .B2(_04229_),
    .X(_04327_));
 sky130_fd_sc_hd__inv_2 _19071_ (.A(\CPU_Dmem_value_a5[12][17] ),
    .Y(_04328_));
 sky130_fd_sc_hd__a2bb2o_4 _19072_ (.A1_N(_04328_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][17] ),
    .B2(_04232_),
    .X(_04329_));
 sky130_fd_sc_hd__or4_4 _19073_ (.A(_04323_),
    .B(_04325_),
    .C(_04327_),
    .D(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__o22a_4 _19074_ (.A1(\CPU_Dmem_value_a5[0][17] ),
    .A2(_04206_),
    .B1(_04321_),
    .B2(_04330_),
    .X(\CPU_dmem_rd_data_a4[17] ));
 sky130_fd_sc_hd__buf_2 _19075_ (.A(_03947_),
    .X(_04331_));
 sky130_fd_sc_hd__inv_2 _19076_ (.A(\CPU_Dmem_value_a5[9][18] ),
    .Y(_04332_));
 sky130_fd_sc_hd__buf_2 _19077_ (.A(_03949_),
    .X(_04333_));
 sky130_fd_sc_hd__buf_2 _19078_ (.A(_03952_),
    .X(_04334_));
 sky130_fd_sc_hd__a2bb2o_4 _19079_ (.A1_N(_04332_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][18] ),
    .B2(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__inv_2 _19080_ (.A(\CPU_Dmem_value_a5[8][18] ),
    .Y(_04336_));
 sky130_fd_sc_hd__buf_2 _19081_ (.A(_03956_),
    .X(_04337_));
 sky130_fd_sc_hd__buf_2 _19082_ (.A(_03959_),
    .X(_04338_));
 sky130_fd_sc_hd__a2bb2o_4 _19083_ (.A1_N(_04336_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][18] ),
    .B2(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__inv_2 _19084_ (.A(\CPU_Dmem_value_a5[2][18] ),
    .Y(_04340_));
 sky130_fd_sc_hd__buf_2 _19085_ (.A(_03963_),
    .X(_04341_));
 sky130_fd_sc_hd__o21ai_4 _19086_ (.A1(_04340_),
    .A2(_04341_),
    .B1(_04299_),
    .Y(_04342_));
 sky130_fd_sc_hd__inv_2 _19087_ (.A(\CPU_Dmem_value_a5[3][18] ),
    .Y(_04343_));
 sky130_fd_sc_hd__buf_2 _19088_ (.A(_03966_),
    .X(_04344_));
 sky130_fd_sc_hd__buf_2 _19089_ (.A(_03969_),
    .X(_04345_));
 sky130_fd_sc_hd__a2bb2o_4 _19090_ (.A1_N(_04343_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][18] ),
    .B2(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__or4_4 _19091_ (.A(_04335_),
    .B(_04339_),
    .C(_04342_),
    .D(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__inv_2 _19092_ (.A(\CPU_Dmem_value_a5[1][18] ),
    .Y(_04348_));
 sky130_fd_sc_hd__a2bb2o_4 _19093_ (.A1_N(_04348_),
    .A2_N(_04245_),
    .B1(\CPU_Dmem_value_a5[4][18] ),
    .B2(_04246_),
    .X(_04349_));
 sky130_fd_sc_hd__inv_2 _19094_ (.A(\CPU_Dmem_value_a5[6][18] ),
    .Y(_04350_));
 sky130_fd_sc_hd__buf_2 _19095_ (.A(_04098_),
    .X(_04351_));
 sky130_fd_sc_hd__a2bb2o_4 _19096_ (.A1_N(_04350_),
    .A2_N(_04249_),
    .B1(\CPU_Dmem_value_a5[11][18] ),
    .B2(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__inv_2 _19097_ (.A(\CPU_Dmem_value_a5[14][18] ),
    .Y(_04353_));
 sky130_fd_sc_hd__buf_2 _19098_ (.A(_04102_),
    .X(_04354_));
 sky130_fd_sc_hd__a2bb2o_4 _19099_ (.A1_N(_04353_),
    .A2_N(_04252_),
    .B1(\CPU_Dmem_value_a5[5][18] ),
    .B2(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__inv_2 _19100_ (.A(\CPU_Dmem_value_a5[12][18] ),
    .Y(_04356_));
 sky130_fd_sc_hd__buf_2 _19101_ (.A(_04106_),
    .X(_04357_));
 sky130_fd_sc_hd__a2bb2o_4 _19102_ (.A1_N(_04356_),
    .A2_N(_04255_),
    .B1(\CPU_Dmem_value_a5[15][18] ),
    .B2(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__or4_4 _19103_ (.A(_04349_),
    .B(_04352_),
    .C(_04355_),
    .D(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__o22a_4 _19104_ (.A1(\CPU_Dmem_value_a5[0][18] ),
    .A2(_04331_),
    .B1(_04347_),
    .B2(_04359_),
    .X(\CPU_dmem_rd_data_a4[18] ));
 sky130_fd_sc_hd__inv_2 _19105_ (.A(\CPU_Dmem_value_a5[9][19] ),
    .Y(_04360_));
 sky130_fd_sc_hd__a2bb2o_4 _19106_ (.A1_N(_04360_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][19] ),
    .B2(_04334_),
    .X(_04361_));
 sky130_fd_sc_hd__inv_2 _19107_ (.A(\CPU_Dmem_value_a5[8][19] ),
    .Y(_04362_));
 sky130_fd_sc_hd__a2bb2o_4 _19108_ (.A1_N(_04362_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][19] ),
    .B2(_04338_),
    .X(_04363_));
 sky130_fd_sc_hd__inv_2 _19109_ (.A(\CPU_Dmem_value_a5[2][19] ),
    .Y(_04364_));
 sky130_fd_sc_hd__o21ai_4 _19110_ (.A1(_04364_),
    .A2(_04341_),
    .B1(_04299_),
    .Y(_04365_));
 sky130_fd_sc_hd__inv_2 _19111_ (.A(\CPU_Dmem_value_a5[3][19] ),
    .Y(_04366_));
 sky130_fd_sc_hd__a2bb2o_4 _19112_ (.A1_N(_04366_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][19] ),
    .B2(_04345_),
    .X(_04367_));
 sky130_fd_sc_hd__or4_4 _19113_ (.A(_04361_),
    .B(_04363_),
    .C(_04365_),
    .D(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__inv_2 _19114_ (.A(\CPU_Dmem_value_a5[1][19] ),
    .Y(_04369_));
 sky130_fd_sc_hd__buf_2 _19115_ (.A(_03973_),
    .X(_04370_));
 sky130_fd_sc_hd__buf_2 _19116_ (.A(_04001_),
    .X(_04371_));
 sky130_fd_sc_hd__a2bb2o_4 _19117_ (.A1_N(_04369_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][19] ),
    .B2(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__inv_2 _19118_ (.A(\CPU_Dmem_value_a5[6][19] ),
    .Y(_04373_));
 sky130_fd_sc_hd__buf_2 _19119_ (.A(_03975_),
    .X(_04374_));
 sky130_fd_sc_hd__a2bb2o_4 _19120_ (.A1_N(_04373_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][19] ),
    .B2(_04351_),
    .X(_04375_));
 sky130_fd_sc_hd__inv_2 _19121_ (.A(\CPU_Dmem_value_a5[14][19] ),
    .Y(_04376_));
 sky130_fd_sc_hd__buf_2 _19122_ (.A(_03980_),
    .X(_04377_));
 sky130_fd_sc_hd__a2bb2o_4 _19123_ (.A1_N(_04376_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][19] ),
    .B2(_04354_),
    .X(_04378_));
 sky130_fd_sc_hd__inv_2 _19124_ (.A(\CPU_Dmem_value_a5[12][19] ),
    .Y(_04379_));
 sky130_fd_sc_hd__buf_2 _19125_ (.A(_03985_),
    .X(_04380_));
 sky130_fd_sc_hd__a2bb2o_4 _19126_ (.A1_N(_04379_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][19] ),
    .B2(_04357_),
    .X(_04381_));
 sky130_fd_sc_hd__or4_4 _19127_ (.A(_04372_),
    .B(_04375_),
    .C(_04378_),
    .D(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__o22a_4 _19128_ (.A1(\CPU_Dmem_value_a5[0][19] ),
    .A2(_04331_),
    .B1(_04368_),
    .B2(_04382_),
    .X(\CPU_dmem_rd_data_a4[19] ));
 sky130_fd_sc_hd__inv_2 _19129_ (.A(\CPU_Dmem_value_a5[9][20] ),
    .Y(_04383_));
 sky130_fd_sc_hd__a2bb2o_4 _19130_ (.A1_N(_04383_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][20] ),
    .B2(_04334_),
    .X(_04384_));
 sky130_fd_sc_hd__inv_2 _19131_ (.A(\CPU_Dmem_value_a5[8][20] ),
    .Y(_04385_));
 sky130_fd_sc_hd__a2bb2o_4 _19132_ (.A1_N(_04385_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][20] ),
    .B2(_04338_),
    .X(_04386_));
 sky130_fd_sc_hd__inv_2 _19133_ (.A(\CPU_Dmem_value_a5[2][20] ),
    .Y(_04387_));
 sky130_fd_sc_hd__o21ai_4 _19134_ (.A1(_04387_),
    .A2(_04341_),
    .B1(_04299_),
    .Y(_04388_));
 sky130_fd_sc_hd__inv_2 _19135_ (.A(\CPU_Dmem_value_a5[3][20] ),
    .Y(_04389_));
 sky130_fd_sc_hd__a2bb2o_4 _19136_ (.A1_N(_04389_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][20] ),
    .B2(_04345_),
    .X(_04390_));
 sky130_fd_sc_hd__or4_4 _19137_ (.A(_04384_),
    .B(_04386_),
    .C(_04388_),
    .D(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__inv_2 _19138_ (.A(\CPU_Dmem_value_a5[1][20] ),
    .Y(_04392_));
 sky130_fd_sc_hd__a2bb2o_4 _19139_ (.A1_N(_04392_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][20] ),
    .B2(_04371_),
    .X(_04393_));
 sky130_fd_sc_hd__inv_2 _19140_ (.A(\CPU_Dmem_value_a5[6][20] ),
    .Y(_04394_));
 sky130_fd_sc_hd__a2bb2o_4 _19141_ (.A1_N(_04394_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][20] ),
    .B2(_04351_),
    .X(_04395_));
 sky130_fd_sc_hd__inv_2 _19142_ (.A(\CPU_Dmem_value_a5[14][20] ),
    .Y(_04396_));
 sky130_fd_sc_hd__a2bb2o_4 _19143_ (.A1_N(_04396_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][20] ),
    .B2(_04354_),
    .X(_04397_));
 sky130_fd_sc_hd__inv_2 _19144_ (.A(\CPU_Dmem_value_a5[12][20] ),
    .Y(_04398_));
 sky130_fd_sc_hd__a2bb2o_4 _19145_ (.A1_N(_04398_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][20] ),
    .B2(_04357_),
    .X(_04399_));
 sky130_fd_sc_hd__or4_4 _19146_ (.A(_04393_),
    .B(_04395_),
    .C(_04397_),
    .D(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__o22a_4 _19147_ (.A1(\CPU_Dmem_value_a5[0][20] ),
    .A2(_04331_),
    .B1(_04391_),
    .B2(_04400_),
    .X(\CPU_dmem_rd_data_a4[20] ));
 sky130_fd_sc_hd__inv_2 _19148_ (.A(\CPU_Dmem_value_a5[9][21] ),
    .Y(_04401_));
 sky130_fd_sc_hd__a2bb2o_4 _19149_ (.A1_N(_04401_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][21] ),
    .B2(_04334_),
    .X(_04402_));
 sky130_fd_sc_hd__inv_2 _19150_ (.A(\CPU_Dmem_value_a5[8][21] ),
    .Y(_04403_));
 sky130_fd_sc_hd__a2bb2o_4 _19151_ (.A1_N(_04403_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][21] ),
    .B2(_04338_),
    .X(_04404_));
 sky130_fd_sc_hd__inv_2 _19152_ (.A(\CPU_Dmem_value_a5[2][21] ),
    .Y(_04405_));
 sky130_fd_sc_hd__o21ai_4 _19153_ (.A1(_04405_),
    .A2(_04341_),
    .B1(_04299_),
    .Y(_04406_));
 sky130_fd_sc_hd__inv_2 _19154_ (.A(\CPU_Dmem_value_a5[3][21] ),
    .Y(_04407_));
 sky130_fd_sc_hd__a2bb2o_4 _19155_ (.A1_N(_04407_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][21] ),
    .B2(_04345_),
    .X(_04408_));
 sky130_fd_sc_hd__or4_4 _19156_ (.A(_04402_),
    .B(_04404_),
    .C(_04406_),
    .D(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__inv_2 _19157_ (.A(\CPU_Dmem_value_a5[1][21] ),
    .Y(_04410_));
 sky130_fd_sc_hd__a2bb2o_4 _19158_ (.A1_N(_04410_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][21] ),
    .B2(_04371_),
    .X(_04411_));
 sky130_fd_sc_hd__inv_2 _19159_ (.A(\CPU_Dmem_value_a5[6][21] ),
    .Y(_04412_));
 sky130_fd_sc_hd__a2bb2o_4 _19160_ (.A1_N(_04412_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][21] ),
    .B2(_04351_),
    .X(_04413_));
 sky130_fd_sc_hd__inv_2 _19161_ (.A(\CPU_Dmem_value_a5[14][21] ),
    .Y(_04414_));
 sky130_fd_sc_hd__a2bb2o_4 _19162_ (.A1_N(_04414_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][21] ),
    .B2(_04354_),
    .X(_04415_));
 sky130_fd_sc_hd__inv_2 _19163_ (.A(\CPU_Dmem_value_a5[12][21] ),
    .Y(_04416_));
 sky130_fd_sc_hd__a2bb2o_4 _19164_ (.A1_N(_04416_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][21] ),
    .B2(_04357_),
    .X(_04417_));
 sky130_fd_sc_hd__or4_4 _19165_ (.A(_04411_),
    .B(_04413_),
    .C(_04415_),
    .D(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__o22a_4 _19166_ (.A1(\CPU_Dmem_value_a5[0][21] ),
    .A2(_04331_),
    .B1(_04409_),
    .B2(_04418_),
    .X(\CPU_dmem_rd_data_a4[21] ));
 sky130_fd_sc_hd__inv_2 _19167_ (.A(\CPU_Dmem_value_a5[9][22] ),
    .Y(_04419_));
 sky130_fd_sc_hd__a2bb2o_4 _19168_ (.A1_N(_04419_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][22] ),
    .B2(_04334_),
    .X(_04420_));
 sky130_fd_sc_hd__inv_2 _19169_ (.A(\CPU_Dmem_value_a5[8][22] ),
    .Y(_04421_));
 sky130_fd_sc_hd__a2bb2o_4 _19170_ (.A1_N(_04421_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][22] ),
    .B2(_04338_),
    .X(_04422_));
 sky130_fd_sc_hd__inv_2 _19171_ (.A(\CPU_Dmem_value_a5[2][22] ),
    .Y(_04423_));
 sky130_fd_sc_hd__buf_2 _19172_ (.A(_04655_),
    .X(_04424_));
 sky130_fd_sc_hd__o21ai_4 _19173_ (.A1(_04423_),
    .A2(_04341_),
    .B1(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__inv_2 _19174_ (.A(\CPU_Dmem_value_a5[3][22] ),
    .Y(_04426_));
 sky130_fd_sc_hd__a2bb2o_4 _19175_ (.A1_N(_04426_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][22] ),
    .B2(_04345_),
    .X(_04427_));
 sky130_fd_sc_hd__or4_4 _19176_ (.A(_04420_),
    .B(_04422_),
    .C(_04425_),
    .D(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__inv_2 _19177_ (.A(\CPU_Dmem_value_a5[1][22] ),
    .Y(_04429_));
 sky130_fd_sc_hd__a2bb2o_4 _19178_ (.A1_N(_04429_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][22] ),
    .B2(_04371_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _19179_ (.A(\CPU_Dmem_value_a5[6][22] ),
    .Y(_04431_));
 sky130_fd_sc_hd__a2bb2o_4 _19180_ (.A1_N(_04431_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][22] ),
    .B2(_04351_),
    .X(_04432_));
 sky130_fd_sc_hd__inv_2 _19181_ (.A(\CPU_Dmem_value_a5[14][22] ),
    .Y(_04433_));
 sky130_fd_sc_hd__a2bb2o_4 _19182_ (.A1_N(_04433_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][22] ),
    .B2(_04354_),
    .X(_04434_));
 sky130_fd_sc_hd__inv_2 _19183_ (.A(\CPU_Dmem_value_a5[12][22] ),
    .Y(_04435_));
 sky130_fd_sc_hd__a2bb2o_4 _19184_ (.A1_N(_04435_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][22] ),
    .B2(_04357_),
    .X(_04436_));
 sky130_fd_sc_hd__or4_4 _19185_ (.A(_04430_),
    .B(_04432_),
    .C(_04434_),
    .D(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__o22a_4 _19186_ (.A1(\CPU_Dmem_value_a5[0][22] ),
    .A2(_04331_),
    .B1(_04428_),
    .B2(_04437_),
    .X(\CPU_dmem_rd_data_a4[22] ));
 sky130_fd_sc_hd__inv_2 _19187_ (.A(\CPU_Dmem_value_a5[9][23] ),
    .Y(_04438_));
 sky130_fd_sc_hd__a2bb2o_4 _19188_ (.A1_N(_04438_),
    .A2_N(_04333_),
    .B1(\CPU_Dmem_value_a5[7][23] ),
    .B2(_04334_),
    .X(_04439_));
 sky130_fd_sc_hd__inv_2 _19189_ (.A(\CPU_Dmem_value_a5[8][23] ),
    .Y(_04440_));
 sky130_fd_sc_hd__a2bb2o_4 _19190_ (.A1_N(_04440_),
    .A2_N(_04337_),
    .B1(\CPU_Dmem_value_a5[13][23] ),
    .B2(_04338_),
    .X(_04441_));
 sky130_fd_sc_hd__inv_2 _19191_ (.A(\CPU_Dmem_value_a5[2][23] ),
    .Y(_04442_));
 sky130_fd_sc_hd__o21ai_4 _19192_ (.A1(_04442_),
    .A2(_04341_),
    .B1(_04424_),
    .Y(_04443_));
 sky130_fd_sc_hd__inv_2 _19193_ (.A(\CPU_Dmem_value_a5[3][23] ),
    .Y(_04444_));
 sky130_fd_sc_hd__a2bb2o_4 _19194_ (.A1_N(_04444_),
    .A2_N(_04344_),
    .B1(\CPU_Dmem_value_a5[10][23] ),
    .B2(_04345_),
    .X(_04445_));
 sky130_fd_sc_hd__or4_4 _19195_ (.A(_04439_),
    .B(_04441_),
    .C(_04443_),
    .D(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__inv_2 _19196_ (.A(\CPU_Dmem_value_a5[1][23] ),
    .Y(_04447_));
 sky130_fd_sc_hd__a2bb2o_4 _19197_ (.A1_N(_04447_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][23] ),
    .B2(_04371_),
    .X(_04448_));
 sky130_fd_sc_hd__inv_2 _19198_ (.A(\CPU_Dmem_value_a5[6][23] ),
    .Y(_04449_));
 sky130_fd_sc_hd__a2bb2o_4 _19199_ (.A1_N(_04449_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][23] ),
    .B2(_04351_),
    .X(_04450_));
 sky130_fd_sc_hd__inv_2 _19200_ (.A(\CPU_Dmem_value_a5[14][23] ),
    .Y(_04451_));
 sky130_fd_sc_hd__a2bb2o_4 _19201_ (.A1_N(_04451_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][23] ),
    .B2(_04354_),
    .X(_04452_));
 sky130_fd_sc_hd__inv_2 _19202_ (.A(\CPU_Dmem_value_a5[12][23] ),
    .Y(_04453_));
 sky130_fd_sc_hd__a2bb2o_4 _19203_ (.A1_N(_04453_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][23] ),
    .B2(_04357_),
    .X(_04454_));
 sky130_fd_sc_hd__or4_4 _19204_ (.A(_04448_),
    .B(_04450_),
    .C(_04452_),
    .D(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__o22a_4 _19205_ (.A1(\CPU_Dmem_value_a5[0][23] ),
    .A2(_04331_),
    .B1(_04446_),
    .B2(_04455_),
    .X(\CPU_dmem_rd_data_a4[23] ));
 sky130_fd_sc_hd__buf_2 _19206_ (.A(_03946_),
    .X(_04456_));
 sky130_fd_sc_hd__inv_2 _19207_ (.A(\CPU_Dmem_value_a5[9][24] ),
    .Y(_04457_));
 sky130_fd_sc_hd__buf_2 _19208_ (.A(_05521_),
    .X(_04458_));
 sky130_fd_sc_hd__buf_2 _19209_ (.A(_03951_),
    .X(_04459_));
 sky130_fd_sc_hd__a2bb2o_4 _19210_ (.A1_N(_04457_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][24] ),
    .B2(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__inv_2 _19211_ (.A(\CPU_Dmem_value_a5[8][24] ),
    .Y(_04461_));
 sky130_fd_sc_hd__buf_2 _19212_ (.A(_05434_),
    .X(_04462_));
 sky130_fd_sc_hd__buf_2 _19213_ (.A(_03958_),
    .X(_04463_));
 sky130_fd_sc_hd__a2bb2o_4 _19214_ (.A1_N(_04461_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][24] ),
    .B2(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__inv_2 _19215_ (.A(\CPU_Dmem_value_a5[2][24] ),
    .Y(_04465_));
 sky130_fd_sc_hd__buf_2 _19216_ (.A(_04895_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_4 _19217_ (.A1(_04465_),
    .A2(_04466_),
    .B1(_04424_),
    .Y(_04467_));
 sky130_fd_sc_hd__inv_2 _19218_ (.A(\CPU_Dmem_value_a5[3][24] ),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_2 _19219_ (.A(_04982_),
    .X(_04469_));
 sky130_fd_sc_hd__buf_2 _19220_ (.A(_03968_),
    .X(_04470_));
 sky130_fd_sc_hd__a2bb2o_4 _19221_ (.A1_N(_04468_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][24] ),
    .B2(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__or4_4 _19222_ (.A(_04460_),
    .B(_04464_),
    .C(_04467_),
    .D(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__inv_2 _19223_ (.A(\CPU_Dmem_value_a5[1][24] ),
    .Y(_04473_));
 sky130_fd_sc_hd__a2bb2o_4 _19224_ (.A1_N(_04473_),
    .A2_N(_04370_),
    .B1(\CPU_Dmem_value_a5[4][24] ),
    .B2(_04371_),
    .X(_04474_));
 sky130_fd_sc_hd__inv_2 _19225_ (.A(\CPU_Dmem_value_a5[6][24] ),
    .Y(_04475_));
 sky130_fd_sc_hd__buf_2 _19226_ (.A(_04098_),
    .X(_04476_));
 sky130_fd_sc_hd__a2bb2o_4 _19227_ (.A1_N(_04475_),
    .A2_N(_04374_),
    .B1(\CPU_Dmem_value_a5[11][24] ),
    .B2(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__inv_2 _19228_ (.A(\CPU_Dmem_value_a5[14][24] ),
    .Y(_04478_));
 sky130_fd_sc_hd__buf_2 _19229_ (.A(_04102_),
    .X(_04479_));
 sky130_fd_sc_hd__a2bb2o_4 _19230_ (.A1_N(_04478_),
    .A2_N(_04377_),
    .B1(\CPU_Dmem_value_a5[5][24] ),
    .B2(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__inv_2 _19231_ (.A(\CPU_Dmem_value_a5[12][24] ),
    .Y(_04481_));
 sky130_fd_sc_hd__buf_2 _19232_ (.A(_04106_),
    .X(_04482_));
 sky130_fd_sc_hd__a2bb2o_4 _19233_ (.A1_N(_04481_),
    .A2_N(_04380_),
    .B1(\CPU_Dmem_value_a5[15][24] ),
    .B2(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__or4_4 _19234_ (.A(_04474_),
    .B(_04477_),
    .C(_04480_),
    .D(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__o22a_4 _19235_ (.A1(\CPU_Dmem_value_a5[0][24] ),
    .A2(_04456_),
    .B1(_04472_),
    .B2(_04484_),
    .X(\CPU_dmem_rd_data_a4[24] ));
 sky130_fd_sc_hd__inv_2 _19236_ (.A(\CPU_Dmem_value_a5[9][25] ),
    .Y(_04485_));
 sky130_fd_sc_hd__a2bb2o_4 _19237_ (.A1_N(_04485_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][25] ),
    .B2(_04459_),
    .X(_04486_));
 sky130_fd_sc_hd__inv_2 _19238_ (.A(\CPU_Dmem_value_a5[8][25] ),
    .Y(_04487_));
 sky130_fd_sc_hd__a2bb2o_4 _19239_ (.A1_N(_04487_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][25] ),
    .B2(_04463_),
    .X(_04488_));
 sky130_fd_sc_hd__inv_2 _19240_ (.A(\CPU_Dmem_value_a5[2][25] ),
    .Y(_04489_));
 sky130_fd_sc_hd__o21ai_4 _19241_ (.A1(_04489_),
    .A2(_04466_),
    .B1(_04424_),
    .Y(_04490_));
 sky130_fd_sc_hd__inv_2 _19242_ (.A(\CPU_Dmem_value_a5[3][25] ),
    .Y(_04491_));
 sky130_fd_sc_hd__a2bb2o_4 _19243_ (.A1_N(_04491_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][25] ),
    .B2(_04470_),
    .X(_04492_));
 sky130_fd_sc_hd__or4_4 _19244_ (.A(_04486_),
    .B(_04488_),
    .C(_04490_),
    .D(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__inv_2 _19245_ (.A(\CPU_Dmem_value_a5[1][25] ),
    .Y(_04494_));
 sky130_fd_sc_hd__buf_2 _19246_ (.A(_04806_),
    .X(_04495_));
 sky130_fd_sc_hd__buf_2 _19247_ (.A(_04001_),
    .X(_04496_));
 sky130_fd_sc_hd__a2bb2o_4 _19248_ (.A1_N(_04494_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][25] ),
    .B2(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__inv_2 _19249_ (.A(\CPU_Dmem_value_a5[6][25] ),
    .Y(_04498_));
 sky130_fd_sc_hd__buf_2 _19250_ (.A(_05239_),
    .X(_04499_));
 sky130_fd_sc_hd__a2bb2o_4 _19251_ (.A1_N(_04498_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][25] ),
    .B2(_04476_),
    .X(_04500_));
 sky130_fd_sc_hd__inv_2 _19252_ (.A(\CPU_Dmem_value_a5[14][25] ),
    .Y(_04501_));
 sky130_fd_sc_hd__buf_2 _19253_ (.A(_05938_),
    .X(_04502_));
 sky130_fd_sc_hd__a2bb2o_4 _19254_ (.A1_N(_04501_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][25] ),
    .B2(_04479_),
    .X(_04503_));
 sky130_fd_sc_hd__inv_2 _19255_ (.A(\CPU_Dmem_value_a5[12][25] ),
    .Y(_04504_));
 sky130_fd_sc_hd__buf_2 _19256_ (.A(_05772_),
    .X(_04505_));
 sky130_fd_sc_hd__a2bb2o_4 _19257_ (.A1_N(_04504_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][25] ),
    .B2(_04482_),
    .X(_04506_));
 sky130_fd_sc_hd__or4_4 _19258_ (.A(_04497_),
    .B(_04500_),
    .C(_04503_),
    .D(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__o22a_4 _19259_ (.A1(\CPU_Dmem_value_a5[0][25] ),
    .A2(_04456_),
    .B1(_04493_),
    .B2(_04507_),
    .X(\CPU_dmem_rd_data_a4[25] ));
 sky130_fd_sc_hd__inv_2 _19260_ (.A(\CPU_Dmem_value_a5[9][26] ),
    .Y(_04508_));
 sky130_fd_sc_hd__a2bb2o_4 _19261_ (.A1_N(_04508_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][26] ),
    .B2(_04459_),
    .X(_04509_));
 sky130_fd_sc_hd__inv_2 _19262_ (.A(\CPU_Dmem_value_a5[8][26] ),
    .Y(_04510_));
 sky130_fd_sc_hd__a2bb2o_4 _19263_ (.A1_N(_04510_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][26] ),
    .B2(_04463_),
    .X(_04511_));
 sky130_fd_sc_hd__inv_2 _19264_ (.A(\CPU_Dmem_value_a5[2][26] ),
    .Y(_04512_));
 sky130_fd_sc_hd__o21ai_4 _19265_ (.A1(_04512_),
    .A2(_04466_),
    .B1(_04424_),
    .Y(_04513_));
 sky130_fd_sc_hd__inv_2 _19266_ (.A(\CPU_Dmem_value_a5[3][26] ),
    .Y(_04514_));
 sky130_fd_sc_hd__a2bb2o_4 _19267_ (.A1_N(_04514_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][26] ),
    .B2(_04470_),
    .X(_04515_));
 sky130_fd_sc_hd__or4_4 _19268_ (.A(_04509_),
    .B(_04511_),
    .C(_04513_),
    .D(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__inv_2 _19269_ (.A(\CPU_Dmem_value_a5[1][26] ),
    .Y(_04517_));
 sky130_fd_sc_hd__a2bb2o_4 _19270_ (.A1_N(_04517_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][26] ),
    .B2(_04496_),
    .X(_04518_));
 sky130_fd_sc_hd__inv_2 _19271_ (.A(\CPU_Dmem_value_a5[6][26] ),
    .Y(_04519_));
 sky130_fd_sc_hd__a2bb2o_4 _19272_ (.A1_N(_04519_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][26] ),
    .B2(_04476_),
    .X(_04520_));
 sky130_fd_sc_hd__inv_2 _19273_ (.A(\CPU_Dmem_value_a5[14][26] ),
    .Y(_04521_));
 sky130_fd_sc_hd__a2bb2o_4 _19274_ (.A1_N(_04521_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][26] ),
    .B2(_04479_),
    .X(_04522_));
 sky130_fd_sc_hd__inv_2 _19275_ (.A(\CPU_Dmem_value_a5[12][26] ),
    .Y(_04523_));
 sky130_fd_sc_hd__a2bb2o_4 _19276_ (.A1_N(_04523_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][26] ),
    .B2(_04482_),
    .X(_04524_));
 sky130_fd_sc_hd__or4_4 _19277_ (.A(_04518_),
    .B(_04520_),
    .C(_04522_),
    .D(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__o22a_4 _19278_ (.A1(\CPU_Dmem_value_a5[0][26] ),
    .A2(_04456_),
    .B1(_04516_),
    .B2(_04525_),
    .X(\CPU_dmem_rd_data_a4[26] ));
 sky130_fd_sc_hd__inv_2 _19279_ (.A(\CPU_Dmem_value_a5[9][27] ),
    .Y(_04526_));
 sky130_fd_sc_hd__a2bb2o_4 _19280_ (.A1_N(_04526_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][27] ),
    .B2(_04459_),
    .X(_04527_));
 sky130_fd_sc_hd__inv_2 _19281_ (.A(\CPU_Dmem_value_a5[8][27] ),
    .Y(_04528_));
 sky130_fd_sc_hd__a2bb2o_4 _19282_ (.A1_N(_04528_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][27] ),
    .B2(_04463_),
    .X(_04529_));
 sky130_fd_sc_hd__inv_2 _19283_ (.A(\CPU_Dmem_value_a5[2][27] ),
    .Y(_04530_));
 sky130_fd_sc_hd__o21ai_4 _19284_ (.A1(_04530_),
    .A2(_04466_),
    .B1(_04424_),
    .Y(_04531_));
 sky130_fd_sc_hd__inv_2 _19285_ (.A(\CPU_Dmem_value_a5[3][27] ),
    .Y(_04532_));
 sky130_fd_sc_hd__a2bb2o_4 _19286_ (.A1_N(_04532_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][27] ),
    .B2(_04470_),
    .X(_04533_));
 sky130_fd_sc_hd__or4_4 _19287_ (.A(_04527_),
    .B(_04529_),
    .C(_04531_),
    .D(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__inv_2 _19288_ (.A(\CPU_Dmem_value_a5[1][27] ),
    .Y(_04535_));
 sky130_fd_sc_hd__a2bb2o_4 _19289_ (.A1_N(_04535_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][27] ),
    .B2(_04496_),
    .X(_04536_));
 sky130_fd_sc_hd__inv_2 _19290_ (.A(\CPU_Dmem_value_a5[6][27] ),
    .Y(_04537_));
 sky130_fd_sc_hd__a2bb2o_4 _19291_ (.A1_N(_04537_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][27] ),
    .B2(_04476_),
    .X(_04538_));
 sky130_fd_sc_hd__inv_2 _19292_ (.A(\CPU_Dmem_value_a5[14][27] ),
    .Y(_04539_));
 sky130_fd_sc_hd__a2bb2o_4 _19293_ (.A1_N(_04539_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][27] ),
    .B2(_04479_),
    .X(_04540_));
 sky130_fd_sc_hd__inv_2 _19294_ (.A(\CPU_Dmem_value_a5[12][27] ),
    .Y(_04541_));
 sky130_fd_sc_hd__a2bb2o_4 _19295_ (.A1_N(_04541_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][27] ),
    .B2(_04482_),
    .X(_04542_));
 sky130_fd_sc_hd__or4_4 _19296_ (.A(_04536_),
    .B(_04538_),
    .C(_04540_),
    .D(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__o22a_4 _19297_ (.A1(\CPU_Dmem_value_a5[0][27] ),
    .A2(_04456_),
    .B1(_04534_),
    .B2(_04543_),
    .X(\CPU_dmem_rd_data_a4[27] ));
 sky130_fd_sc_hd__inv_2 _19298_ (.A(\CPU_Dmem_value_a5[9][28] ),
    .Y(_04544_));
 sky130_fd_sc_hd__a2bb2o_4 _19299_ (.A1_N(_04544_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][28] ),
    .B2(_04459_),
    .X(_04545_));
 sky130_fd_sc_hd__inv_2 _19300_ (.A(\CPU_Dmem_value_a5[8][28] ),
    .Y(_04546_));
 sky130_fd_sc_hd__a2bb2o_4 _19301_ (.A1_N(_04546_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][28] ),
    .B2(_04463_),
    .X(_04547_));
 sky130_fd_sc_hd__inv_2 _19302_ (.A(\CPU_Dmem_value_a5[2][28] ),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ai_4 _19303_ (.A1(_04548_),
    .A2(_04466_),
    .B1(_03945_),
    .Y(_04549_));
 sky130_fd_sc_hd__inv_2 _19304_ (.A(\CPU_Dmem_value_a5[3][28] ),
    .Y(_04550_));
 sky130_fd_sc_hd__a2bb2o_4 _19305_ (.A1_N(_04550_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][28] ),
    .B2(_04470_),
    .X(_04551_));
 sky130_fd_sc_hd__or4_4 _19306_ (.A(_04545_),
    .B(_04547_),
    .C(_04549_),
    .D(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__inv_2 _19307_ (.A(\CPU_Dmem_value_a5[1][28] ),
    .Y(_04553_));
 sky130_fd_sc_hd__a2bb2o_4 _19308_ (.A1_N(_04553_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][28] ),
    .B2(_04496_),
    .X(_04554_));
 sky130_fd_sc_hd__inv_2 _19309_ (.A(\CPU_Dmem_value_a5[6][28] ),
    .Y(_04555_));
 sky130_fd_sc_hd__a2bb2o_4 _19310_ (.A1_N(_04555_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][28] ),
    .B2(_04476_),
    .X(_04556_));
 sky130_fd_sc_hd__inv_2 _19311_ (.A(\CPU_Dmem_value_a5[14][28] ),
    .Y(_04557_));
 sky130_fd_sc_hd__a2bb2o_4 _19312_ (.A1_N(_04557_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][28] ),
    .B2(_04479_),
    .X(_04558_));
 sky130_fd_sc_hd__inv_2 _19313_ (.A(\CPU_Dmem_value_a5[12][28] ),
    .Y(_04559_));
 sky130_fd_sc_hd__a2bb2o_4 _19314_ (.A1_N(_04559_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][28] ),
    .B2(_04482_),
    .X(_04560_));
 sky130_fd_sc_hd__or4_4 _19315_ (.A(_04554_),
    .B(_04556_),
    .C(_04558_),
    .D(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__o22a_4 _19316_ (.A1(\CPU_Dmem_value_a5[0][28] ),
    .A2(_04456_),
    .B1(_04552_),
    .B2(_04561_),
    .X(\CPU_dmem_rd_data_a4[28] ));
 sky130_fd_sc_hd__inv_2 _19317_ (.A(\CPU_Dmem_value_a5[9][29] ),
    .Y(_04562_));
 sky130_fd_sc_hd__a2bb2o_4 _19318_ (.A1_N(_04562_),
    .A2_N(_04458_),
    .B1(\CPU_Dmem_value_a5[7][29] ),
    .B2(_04459_),
    .X(_04563_));
 sky130_fd_sc_hd__inv_2 _19319_ (.A(\CPU_Dmem_value_a5[8][29] ),
    .Y(_04564_));
 sky130_fd_sc_hd__a2bb2o_4 _19320_ (.A1_N(_04564_),
    .A2_N(_04462_),
    .B1(\CPU_Dmem_value_a5[13][29] ),
    .B2(_04463_),
    .X(_04565_));
 sky130_fd_sc_hd__inv_2 _19321_ (.A(\CPU_Dmem_value_a5[2][29] ),
    .Y(_04566_));
 sky130_fd_sc_hd__o21ai_4 _19322_ (.A1(_04566_),
    .A2(_04466_),
    .B1(_03945_),
    .Y(_04567_));
 sky130_fd_sc_hd__inv_2 _19323_ (.A(\CPU_Dmem_value_a5[3][29] ),
    .Y(_04568_));
 sky130_fd_sc_hd__a2bb2o_4 _19324_ (.A1_N(_04568_),
    .A2_N(_04469_),
    .B1(\CPU_Dmem_value_a5[10][29] ),
    .B2(_04470_),
    .X(_04569_));
 sky130_fd_sc_hd__or4_4 _19325_ (.A(_04563_),
    .B(_04565_),
    .C(_04567_),
    .D(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__inv_2 _19326_ (.A(\CPU_Dmem_value_a5[1][29] ),
    .Y(_04571_));
 sky130_fd_sc_hd__a2bb2o_4 _19327_ (.A1_N(_04571_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][29] ),
    .B2(_04496_),
    .X(_04572_));
 sky130_fd_sc_hd__inv_2 _19328_ (.A(\CPU_Dmem_value_a5[6][29] ),
    .Y(_04573_));
 sky130_fd_sc_hd__a2bb2o_4 _19329_ (.A1_N(_04573_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][29] ),
    .B2(_04476_),
    .X(_04574_));
 sky130_fd_sc_hd__inv_2 _19330_ (.A(\CPU_Dmem_value_a5[14][29] ),
    .Y(_04575_));
 sky130_fd_sc_hd__a2bb2o_4 _19331_ (.A1_N(_04575_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][29] ),
    .B2(_04479_),
    .X(_04576_));
 sky130_fd_sc_hd__inv_2 _19332_ (.A(\CPU_Dmem_value_a5[12][29] ),
    .Y(_04577_));
 sky130_fd_sc_hd__a2bb2o_4 _19333_ (.A1_N(_04577_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][29] ),
    .B2(_04482_),
    .X(_04578_));
 sky130_fd_sc_hd__or4_4 _19334_ (.A(_04572_),
    .B(_04574_),
    .C(_04576_),
    .D(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__o22a_4 _19335_ (.A1(\CPU_Dmem_value_a5[0][29] ),
    .A2(_04456_),
    .B1(_04570_),
    .B2(_04579_),
    .X(\CPU_dmem_rd_data_a4[29] ));
 sky130_fd_sc_hd__inv_2 _19336_ (.A(\CPU_Dmem_value_a5[9][30] ),
    .Y(_04580_));
 sky130_fd_sc_hd__a2bb2o_4 _19337_ (.A1_N(_04580_),
    .A2_N(_03949_),
    .B1(\CPU_Dmem_value_a5[7][30] ),
    .B2(_03952_),
    .X(_04581_));
 sky130_fd_sc_hd__inv_2 _19338_ (.A(\CPU_Dmem_value_a5[8][30] ),
    .Y(_04582_));
 sky130_fd_sc_hd__a2bb2o_4 _19339_ (.A1_N(_04582_),
    .A2_N(_03956_),
    .B1(\CPU_Dmem_value_a5[13][30] ),
    .B2(_03959_),
    .X(_04583_));
 sky130_fd_sc_hd__inv_2 _19340_ (.A(\CPU_Dmem_value_a5[2][30] ),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_4 _19341_ (.A1(_04584_),
    .A2(_03963_),
    .B1(_03945_),
    .Y(_04585_));
 sky130_fd_sc_hd__inv_2 _19342_ (.A(\CPU_Dmem_value_a5[3][30] ),
    .Y(_04586_));
 sky130_fd_sc_hd__a2bb2o_4 _19343_ (.A1_N(_04586_),
    .A2_N(_03966_),
    .B1(\CPU_Dmem_value_a5[10][30] ),
    .B2(_03969_),
    .X(_04587_));
 sky130_fd_sc_hd__or4_4 _19344_ (.A(_04581_),
    .B(_04583_),
    .C(_04585_),
    .D(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__inv_2 _19345_ (.A(\CPU_Dmem_value_a5[1][30] ),
    .Y(_04589_));
 sky130_fd_sc_hd__a2bb2o_4 _19346_ (.A1_N(_04589_),
    .A2_N(_04495_),
    .B1(\CPU_Dmem_value_a5[4][30] ),
    .B2(_04496_),
    .X(_04590_));
 sky130_fd_sc_hd__inv_2 _19347_ (.A(\CPU_Dmem_value_a5[6][30] ),
    .Y(_04591_));
 sky130_fd_sc_hd__a2bb2o_4 _19348_ (.A1_N(_04591_),
    .A2_N(_04499_),
    .B1(\CPU_Dmem_value_a5[11][30] ),
    .B2(_04098_),
    .X(_04592_));
 sky130_fd_sc_hd__inv_2 _19349_ (.A(\CPU_Dmem_value_a5[14][30] ),
    .Y(_04593_));
 sky130_fd_sc_hd__a2bb2o_4 _19350_ (.A1_N(_04593_),
    .A2_N(_04502_),
    .B1(\CPU_Dmem_value_a5[5][30] ),
    .B2(_04102_),
    .X(_04594_));
 sky130_fd_sc_hd__inv_2 _19351_ (.A(\CPU_Dmem_value_a5[12][30] ),
    .Y(_04595_));
 sky130_fd_sc_hd__a2bb2o_4 _19352_ (.A1_N(_04595_),
    .A2_N(_04505_),
    .B1(\CPU_Dmem_value_a5[15][30] ),
    .B2(_04106_),
    .X(_04596_));
 sky130_fd_sc_hd__or4_4 _19353_ (.A(_04590_),
    .B(_04592_),
    .C(_04594_),
    .D(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__o22a_4 _19354_ (.A1(\CPU_Dmem_value_a5[0][30] ),
    .A2(_03947_),
    .B1(_04588_),
    .B2(_04597_),
    .X(\CPU_dmem_rd_data_a4[30] ));
 sky130_fd_sc_hd__inv_2 _19355_ (.A(\CPU_Dmem_value_a5[9][31] ),
    .Y(_04598_));
 sky130_fd_sc_hd__a2bb2o_4 _19356_ (.A1_N(_04598_),
    .A2_N(_03949_),
    .B1(\CPU_Dmem_value_a5[7][31] ),
    .B2(_03952_),
    .X(_04599_));
 sky130_fd_sc_hd__inv_2 _19357_ (.A(\CPU_Dmem_value_a5[8][31] ),
    .Y(_04600_));
 sky130_fd_sc_hd__a2bb2o_4 _19358_ (.A1_N(_04600_),
    .A2_N(_03956_),
    .B1(\CPU_Dmem_value_a5[13][31] ),
    .B2(_03959_),
    .X(_04601_));
 sky130_fd_sc_hd__inv_2 _19359_ (.A(\CPU_Dmem_value_a5[2][31] ),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_4 _19360_ (.A1(_04602_),
    .A2(_03963_),
    .B1(_03945_),
    .Y(_04603_));
 sky130_fd_sc_hd__inv_2 _19361_ (.A(\CPU_Dmem_value_a5[3][31] ),
    .Y(_04604_));
 sky130_fd_sc_hd__a2bb2o_4 _19362_ (.A1_N(_04604_),
    .A2_N(_03966_),
    .B1(\CPU_Dmem_value_a5[10][31] ),
    .B2(_03969_),
    .X(_04605_));
 sky130_fd_sc_hd__or4_4 _19363_ (.A(_04599_),
    .B(_04601_),
    .C(_04603_),
    .D(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__inv_2 _19364_ (.A(\CPU_Dmem_value_a5[1][31] ),
    .Y(_04607_));
 sky130_fd_sc_hd__a2bb2o_4 _19365_ (.A1_N(_04607_),
    .A2_N(_03973_),
    .B1(\CPU_Dmem_value_a5[4][31] ),
    .B2(_04001_),
    .X(_04608_));
 sky130_fd_sc_hd__inv_2 _19366_ (.A(\CPU_Dmem_value_a5[6][31] ),
    .Y(_04609_));
 sky130_fd_sc_hd__a2bb2o_4 _19367_ (.A1_N(_04609_),
    .A2_N(_03975_),
    .B1(\CPU_Dmem_value_a5[11][31] ),
    .B2(_04098_),
    .X(_04610_));
 sky130_fd_sc_hd__inv_2 _19368_ (.A(\CPU_Dmem_value_a5[14][31] ),
    .Y(_04611_));
 sky130_fd_sc_hd__a2bb2o_4 _19369_ (.A1_N(_04611_),
    .A2_N(_03980_),
    .B1(\CPU_Dmem_value_a5[5][31] ),
    .B2(_04102_),
    .X(_04612_));
 sky130_fd_sc_hd__inv_2 _19370_ (.A(\CPU_Dmem_value_a5[12][31] ),
    .Y(_04613_));
 sky130_fd_sc_hd__a2bb2o_4 _19371_ (.A1_N(_04613_),
    .A2_N(_03985_),
    .B1(\CPU_Dmem_value_a5[15][31] ),
    .B2(_04106_),
    .X(_04614_));
 sky130_fd_sc_hd__or4_4 _19372_ (.A(_04608_),
    .B(_04610_),
    .C(_04612_),
    .D(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__o22a_4 _19373_ (.A1(\CPU_Dmem_value_a5[0][31] ),
    .A2(_03947_),
    .B1(_04606_),
    .B2(_04615_),
    .X(\CPU_dmem_rd_data_a4[31] ));
 sky130_fd_sc_hd__and2_4 _19374_ (.A(\CPU_inc_pc_a2[0] ),
    .B(\CPU_imm_a2[0] ),
    .X(_04616_));
 sky130_fd_sc_hd__inv_2 _19375_ (.A(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__inv_2 _19376_ (.A(\CPU_inc_pc_a2[1] ),
    .Y(_04618_));
 sky130_fd_sc_hd__inv_2 _19377_ (.A(\CPU_imm_a2[1] ),
    .Y(_04619_));
 sky130_fd_sc_hd__o22a_4 _19378_ (.A1(_04618_),
    .A2(_04619_),
    .B1(\CPU_inc_pc_a2[1] ),
    .B2(\CPU_imm_a2[1] ),
    .X(_04620_));
 sky130_fd_sc_hd__inv_2 _19379_ (.A(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__o22a_4 _19380_ (.A1(_04617_),
    .A2(_04621_),
    .B1(_04616_),
    .B2(_04620_),
    .X(\CPU_br_tgt_pc_a2[1] ));
 sky130_fd_sc_hd__inv_2 _19381_ (.A(\CPU_pc_a2[2] ),
    .Y(_04622_));
 sky130_fd_sc_hd__inv_2 _19382_ (.A(\CPU_imm_a2[2] ),
    .Y(_04623_));
 sky130_fd_sc_hd__and2_4 _19383_ (.A(_04622_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__a21o_4 _19384_ (.A1(\CPU_pc_a2[2] ),
    .A2(\CPU_imm_a2[2] ),
    .B1(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__o22a_4 _19385_ (.A1(_04618_),
    .A2(_04619_),
    .B1(_04617_),
    .B2(_04621_),
    .X(_04626_));
 sky130_fd_sc_hd__a2bb2o_4 _19386_ (.A1_N(_04625_),
    .A2_N(_04626_),
    .B1(_04625_),
    .B2(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__inv_2 _19387_ (.A(_04627_),
    .Y(\CPU_br_tgt_pc_a2[2] ));
 sky130_fd_sc_hd__inv_2 _19388_ (.A(\CPU_pc_a2[3] ),
    .Y(_04628_));
 sky130_fd_sc_hd__inv_2 _19389_ (.A(\CPU_imm_a2[3] ),
    .Y(_04629_));
 sky130_fd_sc_hd__and2_4 _19390_ (.A(_04628_),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__a21o_4 _19391_ (.A1(\CPU_pc_a2[3] ),
    .A2(\CPU_imm_a2[3] ),
    .B1(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__o22a_4 _19392_ (.A1(_04622_),
    .A2(_04623_),
    .B1(_04624_),
    .B2(_04626_),
    .X(_04632_));
 sky130_fd_sc_hd__a2bb2o_4 _19393_ (.A1_N(_04631_),
    .A2_N(_04632_),
    .B1(_04631_),
    .B2(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__inv_2 _19394_ (.A(_04633_),
    .Y(\CPU_br_tgt_pc_a2[3] ));
 sky130_fd_sc_hd__inv_2 _19395_ (.A(\CPU_pc_a2[4] ),
    .Y(_04634_));
 sky130_fd_sc_hd__inv_2 _19396_ (.A(\CPU_imm_a2[4] ),
    .Y(_04635_));
 sky130_fd_sc_hd__a2bb2o_4 _19397_ (.A1_N(_04634_),
    .A2_N(_04635_),
    .B1(_04634_),
    .B2(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__o22a_4 _19398_ (.A1(_04628_),
    .A2(_04629_),
    .B1(_04630_),
    .B2(_04632_),
    .X(_04637_));
 sky130_fd_sc_hd__a2bb2o_4 _19399_ (.A1_N(_04636_),
    .A2_N(_04637_),
    .B1(_04636_),
    .B2(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__inv_2 _19400_ (.A(_04638_),
    .Y(\CPU_br_tgt_pc_a2[4] ));
 sky130_fd_sc_hd__o22a_4 _19401_ (.A1(_04634_),
    .A2(_04635_),
    .B1(_04636_),
    .B2(_04637_),
    .X(_04639_));
 sky130_fd_sc_hd__inv_2 _19402_ (.A(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__inv_2 _19403_ (.A(\CPU_pc_a2[5] ),
    .Y(_04641_));
 sky130_fd_sc_hd__inv_2 _19404_ (.A(\CPU_imm_a2[10] ),
    .Y(_04642_));
 sky130_fd_sc_hd__o22a_4 _19405_ (.A1(_04641_),
    .A2(\CPU_imm_a2[10] ),
    .B1(\CPU_pc_a2[5] ),
    .B2(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a2bb2o_4 _19406_ (.A1_N(_04640_),
    .A2_N(_04643_),
    .B1(_04640_),
    .B2(_04643_),
    .X(\CPU_br_tgt_pc_a2[5] ));
 sky130_fd_sc_hd__o21a_4 _19407_ (.A1(\CPU_inc_pc_a2[0] ),
    .A2(\CPU_imm_a2[0] ),
    .B1(_04617_),
    .X(\CPU_br_tgt_pc_a2[0] ));
 sky130_fd_sc_hd__nor2_4 _19408_ (.A(\CPU_Dmem_value_a5[0][31] ),
    .B(_04657_),
    .Y(_04644_));
 sky130_fd_sc_hd__a211o_4 _19409_ (.A1(_04801_),
    .A2(_04664_),
    .B1(_04888_),
    .C1(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__inv_2 _19410_ (.A(_04645_),
    .Y(_01549_));
 sky130_fd_sc_hd__conb_1 _19411_ (.LO(CPU_is_slt_a1));
 sky130_fd_sc_hd__conb_1 _19412_ (.LO(CPU_is_slti_a1));
 sky130_fd_sc_hd__dfxtp_4 _19413_ (.D(\CPU_Xreg_value_a4[17][0] ),
    .Q(\CPU_Xreg_value_a5[17][0] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19414_ (.D(\CPU_Xreg_value_a4[17][1] ),
    .Q(\CPU_Xreg_value_a5[17][1] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19415_ (.D(\CPU_Xreg_value_a4[17][2] ),
    .Q(\CPU_Xreg_value_a5[17][2] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19416_ (.D(\CPU_Xreg_value_a4[17][3] ),
    .Q(\CPU_Xreg_value_a5[17][3] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19417_ (.D(\CPU_Xreg_value_a4[17][4] ),
    .Q(\CPU_Xreg_value_a5[17][4] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19418_ (.D(\CPU_Xreg_value_a4[17][5] ),
    .Q(\CPU_Xreg_value_a5[17][5] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19419_ (.D(\CPU_Xreg_value_a4[17][6] ),
    .Q(\CPU_Xreg_value_a5[17][6] ),
    .CLK(clknet_8_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19420_ (.D(\CPU_Xreg_value_a4[17][7] ),
    .Q(\CPU_Xreg_value_a5[17][7] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19421_ (.D(\CPU_Xreg_value_a4[17][8] ),
    .Q(\CPU_Xreg_value_a5[17][8] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19422_ (.D(\CPU_Xreg_value_a4[17][9] ),
    .Q(\CPU_Xreg_value_a5[17][9] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19423_ (.D(\CPU_Xreg_value_a4[17][10] ),
    .Q(\CPU_Xreg_value_a5[17][10] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19424_ (.D(\CPU_Xreg_value_a4[17][11] ),
    .Q(\CPU_Xreg_value_a5[17][11] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19425_ (.D(\CPU_Xreg_value_a4[17][12] ),
    .Q(\CPU_Xreg_value_a5[17][12] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19426_ (.D(\CPU_Xreg_value_a4[17][13] ),
    .Q(\CPU_Xreg_value_a5[17][13] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19427_ (.D(\CPU_Xreg_value_a4[17][14] ),
    .Q(\CPU_Xreg_value_a5[17][14] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19428_ (.D(\CPU_Xreg_value_a4[17][15] ),
    .Q(\CPU_Xreg_value_a5[17][15] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19429_ (.D(\CPU_Xreg_value_a4[17][16] ),
    .Q(\CPU_Xreg_value_a5[17][16] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19430_ (.D(\CPU_Xreg_value_a4[17][17] ),
    .Q(\CPU_Xreg_value_a5[17][17] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19431_ (.D(\CPU_Xreg_value_a4[17][18] ),
    .Q(\CPU_Xreg_value_a5[17][18] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19432_ (.D(\CPU_Xreg_value_a4[17][19] ),
    .Q(\CPU_Xreg_value_a5[17][19] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19433_ (.D(\CPU_Xreg_value_a4[17][20] ),
    .Q(\CPU_Xreg_value_a5[17][20] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19434_ (.D(\CPU_Xreg_value_a4[17][21] ),
    .Q(\CPU_Xreg_value_a5[17][21] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19435_ (.D(\CPU_Xreg_value_a4[17][22] ),
    .Q(\CPU_Xreg_value_a5[17][22] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19436_ (.D(\CPU_Xreg_value_a4[17][23] ),
    .Q(\CPU_Xreg_value_a5[17][23] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19437_ (.D(\CPU_Xreg_value_a4[17][24] ),
    .Q(\CPU_Xreg_value_a5[17][24] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19438_ (.D(\CPU_Xreg_value_a4[17][25] ),
    .Q(\CPU_Xreg_value_a5[17][25] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19439_ (.D(\CPU_Xreg_value_a4[17][26] ),
    .Q(\CPU_Xreg_value_a5[17][26] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19440_ (.D(\CPU_Xreg_value_a4[17][27] ),
    .Q(\CPU_Xreg_value_a5[17][27] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19441_ (.D(\CPU_Xreg_value_a4[17][28] ),
    .Q(\CPU_Xreg_value_a5[17][28] ),
    .CLK(clknet_8_167_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19442_ (.D(\CPU_Xreg_value_a4[17][29] ),
    .Q(\CPU_Xreg_value_a5[17][29] ),
    .CLK(clknet_8_167_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19443_ (.D(\CPU_Xreg_value_a4[17][30] ),
    .Q(\CPU_Xreg_value_a5[17][30] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19444_ (.D(\CPU_Xreg_value_a4[17][31] ),
    .Q(\CPU_Xreg_value_a5[17][31] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19445_ (.D(CPU_valid_taken_br_a4),
    .Q(CPU_valid_taken_br_a5),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19446_ (.D(CPU_valid_taken_br_a3),
    .Q(CPU_valid_taken_br_a4),
    .CLK(clknet_8_251_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19447_ (.D(\gen_clkP_CPU_dmem_rd_en_a5.pwr_en ),
    .Q(CPU_valid_load_a5),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19448_ (.D(CPU_valid_load_a3),
    .Q(\gen_clkP_CPU_dmem_rd_en_a5.pwr_en ),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19449_ (.D(CPU_valid_a3),
    .Q(CPU_valid_a4),
    .CLK(clknet_8_246_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19450_ (.D(\CPU_src2_value_a3[0] ),
    .Q(\CPU_dmem_wr_data_a4[0] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19451_ (.D(\CPU_src2_value_a3[1] ),
    .Q(\CPU_dmem_wr_data_a4[1] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19452_ (.D(\CPU_src2_value_a3[2] ),
    .Q(\CPU_dmem_wr_data_a4[2] ),
    .CLK(clknet_8_219_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19453_ (.D(\CPU_src2_value_a3[3] ),
    .Q(\CPU_dmem_wr_data_a4[3] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19454_ (.D(\CPU_src2_value_a3[4] ),
    .Q(\CPU_dmem_wr_data_a4[4] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19455_ (.D(\CPU_src2_value_a3[5] ),
    .Q(\CPU_dmem_wr_data_a4[5] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19456_ (.D(\CPU_src2_value_a3[6] ),
    .Q(\CPU_dmem_wr_data_a4[6] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19457_ (.D(\CPU_src2_value_a3[7] ),
    .Q(\CPU_dmem_wr_data_a4[7] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19458_ (.D(\CPU_src2_value_a3[8] ),
    .Q(\CPU_dmem_wr_data_a4[8] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19459_ (.D(\CPU_src2_value_a3[9] ),
    .Q(\CPU_dmem_wr_data_a4[9] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19460_ (.D(\CPU_src2_value_a3[10] ),
    .Q(\CPU_dmem_wr_data_a4[10] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19461_ (.D(\CPU_src2_value_a3[11] ),
    .Q(\CPU_dmem_wr_data_a4[11] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19462_ (.D(\CPU_src2_value_a3[12] ),
    .Q(\CPU_dmem_wr_data_a4[12] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19463_ (.D(\CPU_src2_value_a3[13] ),
    .Q(\CPU_dmem_wr_data_a4[13] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19464_ (.D(\CPU_src2_value_a3[14] ),
    .Q(\CPU_dmem_wr_data_a4[14] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19465_ (.D(\CPU_src2_value_a3[15] ),
    .Q(\CPU_dmem_wr_data_a4[15] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19466_ (.D(\CPU_src2_value_a3[16] ),
    .Q(\CPU_dmem_wr_data_a4[16] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19467_ (.D(\CPU_src2_value_a3[17] ),
    .Q(\CPU_dmem_wr_data_a4[17] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19468_ (.D(\CPU_src2_value_a3[18] ),
    .Q(\CPU_dmem_wr_data_a4[18] ),
    .CLK(clknet_8_207_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19469_ (.D(\CPU_src2_value_a3[19] ),
    .Q(\CPU_dmem_wr_data_a4[19] ),
    .CLK(clknet_8_219_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19470_ (.D(\CPU_src2_value_a3[20] ),
    .Q(\CPU_dmem_wr_data_a4[20] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19471_ (.D(\CPU_src2_value_a3[21] ),
    .Q(\CPU_dmem_wr_data_a4[21] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19472_ (.D(\CPU_src2_value_a3[22] ),
    .Q(\CPU_dmem_wr_data_a4[22] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19473_ (.D(\CPU_src2_value_a3[23] ),
    .Q(\CPU_dmem_wr_data_a4[23] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19474_ (.D(\CPU_src2_value_a3[24] ),
    .Q(\CPU_dmem_wr_data_a4[24] ),
    .CLK(clknet_8_244_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19475_ (.D(\CPU_src2_value_a3[25] ),
    .Q(\CPU_dmem_wr_data_a4[25] ),
    .CLK(clknet_8_247_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19476_ (.D(\CPU_src2_value_a3[26] ),
    .Q(\CPU_dmem_wr_data_a4[26] ),
    .CLK(clknet_8_247_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19477_ (.D(\CPU_src2_value_a3[27] ),
    .Q(\CPU_dmem_wr_data_a4[27] ),
    .CLK(clknet_8_244_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19478_ (.D(\CPU_src2_value_a3[28] ),
    .Q(\CPU_dmem_wr_data_a4[28] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19479_ (.D(\CPU_src2_value_a3[29] ),
    .Q(\CPU_dmem_wr_data_a4[29] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19480_ (.D(\CPU_src2_value_a3[30] ),
    .Q(\CPU_dmem_wr_data_a4[30] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19481_ (.D(\CPU_src2_value_a3[31] ),
    .Q(\CPU_dmem_wr_data_a4[31] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19482_ (.D(\CPU_src2_value_a2[0] ),
    .Q(\CPU_src2_value_a3[0] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19483_ (.D(\CPU_src2_value_a2[1] ),
    .Q(\CPU_src2_value_a3[1] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19484_ (.D(\CPU_src2_value_a2[2] ),
    .Q(\CPU_src2_value_a3[2] ),
    .CLK(clknet_8_219_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19485_ (.D(\CPU_src2_value_a2[3] ),
    .Q(\CPU_src2_value_a3[3] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19486_ (.D(\CPU_src2_value_a2[4] ),
    .Q(\CPU_src2_value_a3[4] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19487_ (.D(\CPU_src2_value_a2[5] ),
    .Q(\CPU_src2_value_a3[5] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19488_ (.D(\CPU_src2_value_a2[6] ),
    .Q(\CPU_src2_value_a3[6] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19489_ (.D(\CPU_src2_value_a2[7] ),
    .Q(\CPU_src2_value_a3[7] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19490_ (.D(\CPU_src2_value_a2[8] ),
    .Q(\CPU_src2_value_a3[8] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19491_ (.D(\CPU_src2_value_a2[9] ),
    .Q(\CPU_src2_value_a3[9] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19492_ (.D(\CPU_src2_value_a2[10] ),
    .Q(\CPU_src2_value_a3[10] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19493_ (.D(\CPU_src2_value_a2[11] ),
    .Q(\CPU_src2_value_a3[11] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19494_ (.D(\CPU_src2_value_a2[12] ),
    .Q(\CPU_src2_value_a3[12] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19495_ (.D(\CPU_src2_value_a2[13] ),
    .Q(\CPU_src2_value_a3[13] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19496_ (.D(\CPU_src2_value_a2[14] ),
    .Q(\CPU_src2_value_a3[14] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19497_ (.D(\CPU_src2_value_a2[15] ),
    .Q(\CPU_src2_value_a3[15] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19498_ (.D(\CPU_src2_value_a2[16] ),
    .Q(\CPU_src2_value_a3[16] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19499_ (.D(\CPU_src2_value_a2[17] ),
    .Q(\CPU_src2_value_a3[17] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19500_ (.D(\CPU_src2_value_a2[18] ),
    .Q(\CPU_src2_value_a3[18] ),
    .CLK(clknet_8_206_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19501_ (.D(\CPU_src2_value_a2[19] ),
    .Q(\CPU_src2_value_a3[19] ),
    .CLK(clknet_8_207_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19502_ (.D(\CPU_src2_value_a2[20] ),
    .Q(\CPU_src2_value_a3[20] ),
    .CLK(clknet_8_207_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19503_ (.D(\CPU_src2_value_a2[21] ),
    .Q(\CPU_src2_value_a3[21] ),
    .CLK(clknet_8_207_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19504_ (.D(\CPU_src2_value_a2[22] ),
    .Q(\CPU_src2_value_a3[22] ),
    .CLK(clknet_8_229_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19505_ (.D(\CPU_src2_value_a2[23] ),
    .Q(\CPU_src2_value_a3[23] ),
    .CLK(clknet_8_229_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19506_ (.D(\CPU_src2_value_a2[24] ),
    .Q(\CPU_src2_value_a3[24] ),
    .CLK(clknet_8_231_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19507_ (.D(\CPU_src2_value_a2[25] ),
    .Q(\CPU_src2_value_a3[25] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19508_ (.D(\CPU_src2_value_a2[26] ),
    .Q(\CPU_src2_value_a3[26] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19509_ (.D(\CPU_src2_value_a2[27] ),
    .Q(\CPU_src2_value_a3[27] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19510_ (.D(\CPU_src2_value_a2[28] ),
    .Q(\CPU_src2_value_a3[28] ),
    .CLK(clknet_8_242_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19511_ (.D(\CPU_src2_value_a2[29] ),
    .Q(\CPU_src2_value_a3[29] ),
    .CLK(clknet_8_243_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19512_ (.D(\CPU_src2_value_a2[30] ),
    .Q(\CPU_src2_value_a3[30] ),
    .CLK(clknet_8_218_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19513_ (.D(\CPU_src2_value_a2[31] ),
    .Q(\CPU_src2_value_a3[31] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19514_ (.D(\CPU_src1_value_a2[0] ),
    .Q(\CPU_src1_value_a3[0] ),
    .CLK(clknet_8_218_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19515_ (.D(\CPU_src1_value_a2[1] ),
    .Q(\CPU_src1_value_a3[1] ),
    .CLK(clknet_8_218_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19516_ (.D(\CPU_src1_value_a2[2] ),
    .Q(\CPU_src1_value_a3[2] ),
    .CLK(clknet_8_219_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19517_ (.D(\CPU_src1_value_a2[3] ),
    .Q(\CPU_src1_value_a3[3] ),
    .CLK(clknet_8_217_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19518_ (.D(\CPU_src1_value_a2[4] ),
    .Q(\CPU_src1_value_a3[4] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19519_ (.D(\CPU_src1_value_a2[5] ),
    .Q(\CPU_src1_value_a3[5] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19520_ (.D(\CPU_src1_value_a2[6] ),
    .Q(\CPU_src1_value_a3[6] ),
    .CLK(clknet_8_218_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19521_ (.D(\CPU_src1_value_a2[7] ),
    .Q(\CPU_src1_value_a3[7] ),
    .CLK(clknet_8_216_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19522_ (.D(\CPU_src1_value_a2[8] ),
    .Q(\CPU_src1_value_a3[8] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19523_ (.D(\CPU_src1_value_a2[9] ),
    .Q(\CPU_src1_value_a3[9] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19524_ (.D(\CPU_src1_value_a2[10] ),
    .Q(\CPU_src1_value_a3[10] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19525_ (.D(\CPU_src1_value_a2[11] ),
    .Q(\CPU_src1_value_a3[11] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19526_ (.D(\CPU_src1_value_a2[12] ),
    .Q(\CPU_src1_value_a3[12] ),
    .CLK(clknet_8_204_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19527_ (.D(\CPU_src1_value_a2[13] ),
    .Q(\CPU_src1_value_a3[13] ),
    .CLK(clknet_8_205_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19528_ (.D(\CPU_src1_value_a2[14] ),
    .Q(\CPU_src1_value_a3[14] ),
    .CLK(clknet_8_205_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19529_ (.D(\CPU_src1_value_a2[15] ),
    .Q(\CPU_src1_value_a3[15] ),
    .CLK(clknet_8_205_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19530_ (.D(\CPU_src1_value_a2[16] ),
    .Q(\CPU_src1_value_a3[16] ),
    .CLK(clknet_8_205_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19531_ (.D(\CPU_src1_value_a2[17] ),
    .Q(\CPU_src1_value_a3[17] ),
    .CLK(clknet_8_205_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19532_ (.D(\CPU_src1_value_a2[18] ),
    .Q(\CPU_src1_value_a3[18] ),
    .CLK(clknet_8_229_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19533_ (.D(\CPU_src1_value_a2[19] ),
    .Q(\CPU_src1_value_a3[19] ),
    .CLK(clknet_8_229_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19534_ (.D(\CPU_src1_value_a2[20] ),
    .Q(\CPU_src1_value_a3[20] ),
    .CLK(clknet_8_228_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19535_ (.D(\CPU_src1_value_a2[21] ),
    .Q(\CPU_src1_value_a3[21] ),
    .CLK(clknet_8_228_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19536_ (.D(\CPU_src1_value_a2[22] ),
    .Q(\CPU_src1_value_a3[22] ),
    .CLK(clknet_8_228_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19537_ (.D(\CPU_src1_value_a2[23] ),
    .Q(\CPU_src1_value_a3[23] ),
    .CLK(clknet_8_228_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19538_ (.D(\CPU_src1_value_a2[24] ),
    .Q(\CPU_src1_value_a3[24] ),
    .CLK(clknet_8_231_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19539_ (.D(\CPU_src1_value_a2[25] ),
    .Q(\CPU_src1_value_a3[25] ),
    .CLK(clknet_8_231_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19540_ (.D(\CPU_src1_value_a2[26] ),
    .Q(\CPU_src1_value_a3[26] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19541_ (.D(\CPU_src1_value_a2[27] ),
    .Q(\CPU_src1_value_a3[27] ),
    .CLK(clknet_8_248_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19542_ (.D(\CPU_src1_value_a2[28] ),
    .Q(\CPU_src1_value_a3[28] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19543_ (.D(\CPU_src1_value_a2[29] ),
    .Q(\CPU_src1_value_a3[29] ),
    .CLK(clknet_8_242_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19544_ (.D(\CPU_src1_value_a2[30] ),
    .Q(\CPU_src1_value_a3[30] ),
    .CLK(clknet_8_244_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19545_ (.D(\CPU_src1_value_a2[31] ),
    .Q(\CPU_src1_value_a3[31] ),
    .CLK(clknet_8_244_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19546_ (.D(\CPU_imem_rd_data_a1[20] ),
    .Q(\CPU_rf_rd_index2_a2[0] ),
    .CLK(clknet_8_248_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19547_ (.D(\CPU_imem_rd_data_a1[21] ),
    .Q(\CPU_rf_rd_index2_a2[1] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19548_ (.D(\CPU_imem_rd_data_a1[22] ),
    .Q(\CPU_rf_rd_index2_a2[2] ),
    .CLK(clknet_8_248_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19549_ (.D(\CPU_imem_rd_data_a1[23] ),
    .Q(\CPU_rf_rd_index2_a2[3] ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19550_ (.D(\CPU_imem_rd_data_a1[24] ),
    .Q(\CPU_rf_rd_index2_a2[4] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19551_ (.D(\CPU_imem_rd_data_a1[15] ),
    .Q(\CPU_rf_rd_index1_a2[0] ),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19552_ (.D(\CPU_imem_rd_data_a1[16] ),
    .Q(\CPU_rf_rd_index1_a2[1] ),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19553_ (.D(\CPU_imem_rd_data_a1[17] ),
    .Q(\CPU_rf_rd_index1_a2[2] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19554_ (.D(\CPU_imem_rd_data_a1[18] ),
    .Q(\CPU_rf_rd_index1_a2[3] ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19555_ (.D(\CPU_result_a3[2] ),
    .Q(\CPU_dmem_addr_a4[0] ),
    .CLK(clknet_8_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19556_ (.D(\CPU_result_a3[3] ),
    .Q(\CPU_dmem_addr_a4[1] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19557_ (.D(\CPU_result_a3[4] ),
    .Q(\CPU_dmem_addr_a4[2] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19558_ (.D(\CPU_result_a3[5] ),
    .Q(\CPU_dmem_addr_a4[3] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19559_ (.D(CPU_reset_a3),
    .Q(CPU_reset_a4),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19560_ (.D(CPU_reset_a2),
    .Q(CPU_reset_a3),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19561_ (.D(CPU_reset_a1),
    .Q(CPU_reset_a2),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19562_ (.D(reset),
    .Q(CPU_reset_a1),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19563_ (.D(\gen_clkP_CPU_rd_valid_a3.pwr_en ),
    .Q(\gen_clkP_CPU_rd_valid_a4.pwr_en ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19564_ (.D(\gen_clkP_CPU_rd_valid_a2.pwr_en ),
    .Q(\gen_clkP_CPU_rd_valid_a3.pwr_en ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19565_ (.D(\CPU_rd_a4[0] ),
    .Q(\CPU_rd_a5[0] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19566_ (.D(\CPU_rd_a4[1] ),
    .Q(\CPU_rd_a5[1] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19567_ (.D(\CPU_rd_a4[2] ),
    .Q(\CPU_rd_a5[2] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19568_ (.D(\CPU_rd_a4[3] ),
    .Q(\CPU_rd_a5[3] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19569_ (.D(\CPU_rd_a4[4] ),
    .Q(\CPU_rd_a5[4] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19570_ (.D(\CPU_rd_a3[0] ),
    .Q(\CPU_rd_a4[0] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19571_ (.D(\CPU_rd_a3[1] ),
    .Q(\CPU_rd_a4[1] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19572_ (.D(\CPU_rd_a3[2] ),
    .Q(\CPU_rd_a4[2] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19573_ (.D(\CPU_rd_a3[3] ),
    .Q(\CPU_rd_a4[3] ),
    .CLK(clknet_8_230_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19574_ (.D(\CPU_rd_a3[4] ),
    .Q(\CPU_rd_a4[4] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19575_ (.D(\CPU_rd_a2[0] ),
    .Q(\CPU_rd_a3[0] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19576_ (.D(\CPU_rd_a2[1] ),
    .Q(\CPU_rd_a3[1] ),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19577_ (.D(\CPU_rd_a2[2] ),
    .Q(\CPU_rd_a3[2] ),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19578_ (.D(\CPU_rd_a2[3] ),
    .Q(\CPU_rd_a3[3] ),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19579_ (.D(\CPU_rd_a2[4] ),
    .Q(\CPU_rd_a3[4] ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19580_ (.D(\CPU_imem_rd_data_a1[7] ),
    .Q(\CPU_rd_a2[0] ),
    .CLK(clknet_8_237_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19581_ (.D(\CPU_imem_rd_data_a1[8] ),
    .Q(\CPU_rd_a2[1] ),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19582_ (.D(\CPU_imem_rd_data_a1[9] ),
    .Q(\CPU_rd_a2[2] ),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19583_ (.D(\CPU_imem_rd_data_a1[10] ),
    .Q(\CPU_rd_a2[3] ),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19584_ (.D(\CPU_imem_rd_data_a1[11] ),
    .Q(\CPU_rd_a2[4] ),
    .CLK(clknet_8_236_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19585_ (.D(\CPU_imem_rd_addr_a1[0] ),
    .Q(\CPU_pc_a2[2] ),
    .CLK(clknet_8_252_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19586_ (.D(\CPU_imem_rd_addr_a1[1] ),
    .Q(\CPU_pc_a2[3] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19587_ (.D(\CPU_imem_rd_addr_a1[2] ),
    .Q(\CPU_pc_a2[4] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19588_ (.D(\CPU_imem_rd_addr_a1[3] ),
    .Q(\CPU_pc_a2[5] ),
    .CLK(clknet_8_251_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19589_ (.D(CPU_is_slti_a2),
    .Q(CPU_is_slti_a3),
    .CLK(clknet_8_241_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19590_ (.D(CPU_is_slti_a1),
    .Q(CPU_is_slti_a2),
    .CLK(clknet_8_241_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19591_ (.D(CPU_is_slt_a2),
    .Q(CPU_is_slt_a3),
    .CLK(clknet_8_246_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19592_ (.D(CPU_is_slt_a1),
    .Q(CPU_is_slt_a2),
    .CLK(clknet_8_246_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19593_ (.D(CPU_is_s_instr_a3),
    .Q(CPU_is_s_instr_a4),
    .CLK(clknet_8_247_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19594_ (.D(CPU_is_s_instr_a2),
    .Q(CPU_is_s_instr_a3),
    .CLK(clknet_8_241_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19595_ (.D(CPU_is_s_instr_a1),
    .Q(CPU_is_s_instr_a2),
    .CLK(clknet_8_240_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19596_ (.D(CPU_is_load_a2),
    .Q(CPU_is_load_a3),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19597_ (.D(CPU_is_load_a1),
    .Q(CPU_is_load_a2),
    .CLK(clknet_8_238_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19598_ (.D(CPU_is_bltu_a2),
    .Q(CPU_is_bltu_a3),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19599_ (.D(CPU_is_bltu_a1),
    .Q(CPU_is_bltu_a2),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19600_ (.D(CPU_is_blt_a2),
    .Q(CPU_is_blt_a3),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19601_ (.D(CPU_is_blt_a1),
    .Q(CPU_is_blt_a2),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19602_ (.D(CPU_is_addi_a2),
    .Q(CPU_is_addi_a3),
    .CLK(clknet_8_240_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19603_ (.D(CPU_is_addi_a1),
    .Q(CPU_is_addi_a2),
    .CLK(clknet_8_243_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19604_ (.D(CPU_is_add_a2),
    .Q(CPU_is_add_a3),
    .CLK(clknet_8_240_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19605_ (.D(CPU_is_add_a1),
    .Q(CPU_is_add_a2),
    .CLK(clknet_8_243_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19606_ (.D(\CPU_inc_pc_a2[0] ),
    .Q(\CPU_inc_pc_a3[0] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19607_ (.D(\CPU_inc_pc_a2[1] ),
    .Q(\CPU_inc_pc_a3[1] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19608_ (.D(\CPU_inc_pc_a2[2] ),
    .Q(\CPU_inc_pc_a3[2] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19609_ (.D(\CPU_inc_pc_a2[3] ),
    .Q(\CPU_inc_pc_a3[3] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19610_ (.D(\CPU_inc_pc_a2[4] ),
    .Q(\CPU_inc_pc_a3[4] ),
    .CLK(clknet_8_251_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19611_ (.D(\CPU_inc_pc_a2[5] ),
    .Q(\CPU_inc_pc_a3[5] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19612_ (.D(\CPU_inc_pc_a1[0] ),
    .Q(\CPU_inc_pc_a2[0] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19613_ (.D(\CPU_inc_pc_a1[1] ),
    .Q(\CPU_inc_pc_a2[1] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19614_ (.D(\CPU_inc_pc_a1[2] ),
    .Q(\CPU_inc_pc_a2[2] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19615_ (.D(\CPU_inc_pc_a1[3] ),
    .Q(\CPU_inc_pc_a2[3] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19616_ (.D(\CPU_inc_pc_a1[4] ),
    .Q(\CPU_inc_pc_a2[4] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19617_ (.D(\CPU_inc_pc_a1[5] ),
    .Q(\CPU_inc_pc_a2[5] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19618_ (.D(\CPU_imm_a2[0] ),
    .Q(\CPU_imm_a3[0] ),
    .CLK(clknet_8_247_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19619_ (.D(\CPU_imm_a2[1] ),
    .Q(\CPU_imm_a3[1] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19620_ (.D(\CPU_imm_a2[2] ),
    .Q(\CPU_imm_a3[2] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19621_ (.D(\CPU_imm_a2[3] ),
    .Q(\CPU_imm_a3[3] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19622_ (.D(\CPU_imm_a2[4] ),
    .Q(\CPU_imm_a3[4] ),
    .CLK(clknet_8_243_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19623_ (.D(\CPU_imm_a2[11] ),
    .Q(\CPU_imm_a3[11] ),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19624_ (.D(\CPU_imm_a2[10] ),
    .Q(\CPU_imm_a3[10] ),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19625_ (.D(\CPU_imm_a1[0] ),
    .Q(\CPU_imm_a2[0] ),
    .CLK(clknet_8_242_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19626_ (.D(\CPU_imm_a1[1] ),
    .Q(\CPU_imm_a2[1] ),
    .CLK(clknet_8_248_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19627_ (.D(\CPU_imm_a1[2] ),
    .Q(\CPU_imm_a2[2] ),
    .CLK(clknet_8_252_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19628_ (.D(\CPU_imm_a1[3] ),
    .Q(\CPU_imm_a2[3] ),
    .CLK(clknet_8_252_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19629_ (.D(\CPU_imm_a1[4] ),
    .Q(\CPU_imm_a2[4] ),
    .CLK(clknet_8_252_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19630_ (.D(\CPU_imm_a1[11] ),
    .Q(\CPU_imm_a2[11] ),
    .CLK(clknet_8_248_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19631_ (.D(\CPU_imm_a1[10] ),
    .Q(\CPU_imm_a2[10] ),
    .CLK(clknet_8_249_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19632_ (.D(\CPU_dmem_rd_data_a4[0] ),
    .Q(\CPU_dmem_rd_data_a5[0] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19633_ (.D(\CPU_dmem_rd_data_a4[1] ),
    .Q(\CPU_dmem_rd_data_a5[1] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19634_ (.D(\CPU_dmem_rd_data_a4[2] ),
    .Q(\CPU_dmem_rd_data_a5[2] ),
    .CLK(clknet_8_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19635_ (.D(\CPU_dmem_rd_data_a4[3] ),
    .Q(\CPU_dmem_rd_data_a5[3] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19636_ (.D(\CPU_dmem_rd_data_a4[4] ),
    .Q(\CPU_dmem_rd_data_a5[4] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19637_ (.D(\CPU_dmem_rd_data_a4[5] ),
    .Q(\CPU_dmem_rd_data_a5[5] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19638_ (.D(\CPU_dmem_rd_data_a4[6] ),
    .Q(\CPU_dmem_rd_data_a5[6] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19639_ (.D(\CPU_dmem_rd_data_a4[7] ),
    .Q(\CPU_dmem_rd_data_a5[7] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19640_ (.D(\CPU_dmem_rd_data_a4[8] ),
    .Q(\CPU_dmem_rd_data_a5[8] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19641_ (.D(\CPU_dmem_rd_data_a4[9] ),
    .Q(\CPU_dmem_rd_data_a5[9] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19642_ (.D(\CPU_dmem_rd_data_a4[10] ),
    .Q(\CPU_dmem_rd_data_a5[10] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19643_ (.D(\CPU_dmem_rd_data_a4[11] ),
    .Q(\CPU_dmem_rd_data_a5[11] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19644_ (.D(\CPU_dmem_rd_data_a4[12] ),
    .Q(\CPU_dmem_rd_data_a5[12] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19645_ (.D(\CPU_dmem_rd_data_a4[13] ),
    .Q(\CPU_dmem_rd_data_a5[13] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19646_ (.D(\CPU_dmem_rd_data_a4[14] ),
    .Q(\CPU_dmem_rd_data_a5[14] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19647_ (.D(\CPU_dmem_rd_data_a4[15] ),
    .Q(\CPU_dmem_rd_data_a5[15] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19648_ (.D(\CPU_dmem_rd_data_a4[16] ),
    .Q(\CPU_dmem_rd_data_a5[16] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19649_ (.D(\CPU_dmem_rd_data_a4[17] ),
    .Q(\CPU_dmem_rd_data_a5[17] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19650_ (.D(\CPU_dmem_rd_data_a4[18] ),
    .Q(\CPU_dmem_rd_data_a5[18] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19651_ (.D(\CPU_dmem_rd_data_a4[19] ),
    .Q(\CPU_dmem_rd_data_a5[19] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19652_ (.D(\CPU_dmem_rd_data_a4[20] ),
    .Q(\CPU_dmem_rd_data_a5[20] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19653_ (.D(\CPU_dmem_rd_data_a4[21] ),
    .Q(\CPU_dmem_rd_data_a5[21] ),
    .CLK(clknet_8_204_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19654_ (.D(\CPU_dmem_rd_data_a4[22] ),
    .Q(\CPU_dmem_rd_data_a5[22] ),
    .CLK(clknet_8_204_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19655_ (.D(\CPU_dmem_rd_data_a4[23] ),
    .Q(\CPU_dmem_rd_data_a5[23] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19656_ (.D(\CPU_dmem_rd_data_a4[24] ),
    .Q(\CPU_dmem_rd_data_a5[24] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19657_ (.D(\CPU_dmem_rd_data_a4[25] ),
    .Q(\CPU_dmem_rd_data_a5[25] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19658_ (.D(\CPU_dmem_rd_data_a4[26] ),
    .Q(\CPU_dmem_rd_data_a5[26] ),
    .CLK(clknet_8_244_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19659_ (.D(\CPU_dmem_rd_data_a4[27] ),
    .Q(\CPU_dmem_rd_data_a5[27] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19660_ (.D(\CPU_dmem_rd_data_a4[28] ),
    .Q(\CPU_dmem_rd_data_a5[28] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19661_ (.D(\CPU_dmem_rd_data_a4[29] ),
    .Q(\CPU_dmem_rd_data_a5[29] ),
    .CLK(clknet_8_245_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19662_ (.D(\CPU_dmem_rd_data_a4[30] ),
    .Q(\CPU_dmem_rd_data_a5[30] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19663_ (.D(\CPU_dmem_rd_data_a4[31] ),
    .Q(\CPU_dmem_rd_data_a5[31] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19664_ (.D(\CPU_br_tgt_pc_a2[0] ),
    .Q(\CPU_br_tgt_pc_a3[0] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19665_ (.D(\CPU_br_tgt_pc_a2[1] ),
    .Q(\CPU_br_tgt_pc_a3[1] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19666_ (.D(\CPU_br_tgt_pc_a2[2] ),
    .Q(\CPU_br_tgt_pc_a3[2] ),
    .CLK(clknet_8_252_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19667_ (.D(\CPU_br_tgt_pc_a2[3] ),
    .Q(\CPU_br_tgt_pc_a3[3] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19668_ (.D(\CPU_br_tgt_pc_a2[4] ),
    .Q(\CPU_br_tgt_pc_a3[4] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19669_ (.D(\CPU_br_tgt_pc_a2[5] ),
    .Q(\CPU_br_tgt_pc_a3[5] ),
    .CLK(clknet_8_251_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19670_ (.D(_00000_),
    .Q(out[0]),
    .CLK(clknet_8_239_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19671_ (.D(_00001_),
    .Q(out[1]),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19672_ (.D(_00002_),
    .Q(out[2]),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19673_ (.D(_00003_),
    .Q(out[3]),
    .CLK(clknet_opt_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19674_ (.D(_00004_),
    .Q(out[4]),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19675_ (.D(_00005_),
    .Q(out[5]),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19676_ (.D(_00006_),
    .Q(out[6]),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19677_ (.D(_00007_),
    .Q(out[7]),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19678_ (.D(_00008_),
    .Q(\CPU_imem_rd_addr_a1[0] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19679_ (.D(_00009_),
    .Q(\CPU_imem_rd_addr_a1[1] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19680_ (.D(_00010_),
    .Q(\CPU_imem_rd_addr_a1[2] ),
    .CLK(clknet_8_254_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19681_ (.D(_00011_),
    .Q(\CPU_imem_rd_addr_a1[3] ),
    .CLK(clknet_8_250_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19682_ (.D(_00012_),
    .Q(\CPU_inc_pc_a1[0] ),
    .CLK(clknet_8_255_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19683_ (.D(_00013_),
    .Q(\CPU_inc_pc_a1[1] ),
    .CLK(clknet_8_253_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19684_ (.D(_00014_),
    .Q(\CPU_Xreg_value_a4[31][0] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19685_ (.D(_00015_),
    .Q(\CPU_Xreg_value_a4[31][1] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19686_ (.D(_00016_),
    .Q(\CPU_Xreg_value_a4[31][2] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19687_ (.D(_00017_),
    .Q(\CPU_Xreg_value_a4[31][3] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19688_ (.D(_00018_),
    .Q(\CPU_Xreg_value_a4[31][4] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19689_ (.D(_00019_),
    .Q(\CPU_Xreg_value_a4[31][5] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19690_ (.D(_00020_),
    .Q(\CPU_Xreg_value_a4[31][6] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19691_ (.D(_00021_),
    .Q(\CPU_Xreg_value_a4[31][7] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19692_ (.D(_00022_),
    .Q(\CPU_Xreg_value_a4[31][8] ),
    .CLK(clknet_8_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19693_ (.D(_00023_),
    .Q(\CPU_Xreg_value_a4[31][9] ),
    .CLK(clknet_8_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19694_ (.D(_00024_),
    .Q(\CPU_Xreg_value_a4[31][10] ),
    .CLK(clknet_8_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19695_ (.D(_00025_),
    .Q(\CPU_Xreg_value_a4[31][11] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19696_ (.D(_00026_),
    .Q(\CPU_Xreg_value_a4[31][12] ),
    .CLK(clknet_8_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19697_ (.D(_00027_),
    .Q(\CPU_Xreg_value_a4[31][13] ),
    .CLK(clknet_8_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19698_ (.D(_00028_),
    .Q(\CPU_Xreg_value_a4[31][14] ),
    .CLK(clknet_8_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19699_ (.D(_00029_),
    .Q(\CPU_Xreg_value_a4[31][15] ),
    .CLK(clknet_8_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19700_ (.D(_00030_),
    .Q(\CPU_Xreg_value_a4[31][16] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19701_ (.D(_00031_),
    .Q(\CPU_Xreg_value_a4[31][17] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19702_ (.D(_00032_),
    .Q(\CPU_Xreg_value_a4[31][18] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19703_ (.D(_00033_),
    .Q(\CPU_Xreg_value_a4[31][19] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19704_ (.D(_00034_),
    .Q(\CPU_Xreg_value_a4[31][20] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19705_ (.D(_00035_),
    .Q(\CPU_Xreg_value_a4[31][21] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19706_ (.D(_00036_),
    .Q(\CPU_Xreg_value_a4[31][22] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19707_ (.D(_00037_),
    .Q(\CPU_Xreg_value_a4[31][23] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19708_ (.D(_00038_),
    .Q(\CPU_Xreg_value_a4[31][24] ),
    .CLK(clknet_8_167_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19709_ (.D(_00039_),
    .Q(\CPU_Xreg_value_a4[31][25] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19710_ (.D(_00040_),
    .Q(\CPU_Xreg_value_a4[31][26] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19711_ (.D(_00041_),
    .Q(\CPU_Xreg_value_a4[31][27] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19712_ (.D(_00042_),
    .Q(\CPU_Xreg_value_a4[31][28] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19713_ (.D(_00043_),
    .Q(\CPU_Xreg_value_a4[31][29] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19714_ (.D(_00044_),
    .Q(\CPU_Xreg_value_a4[31][30] ),
    .CLK(clknet_8_167_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19715_ (.D(_00045_),
    .Q(\CPU_Xreg_value_a4[31][31] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19716_ (.D(_00046_),
    .Q(\CPU_Xreg_value_a4[30][0] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19717_ (.D(_00047_),
    .Q(\CPU_Xreg_value_a4[30][1] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19718_ (.D(_00048_),
    .Q(\CPU_Xreg_value_a4[30][2] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19719_ (.D(_00049_),
    .Q(\CPU_Xreg_value_a4[30][3] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19720_ (.D(_00050_),
    .Q(\CPU_Xreg_value_a4[30][4] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19721_ (.D(_00051_),
    .Q(\CPU_Xreg_value_a4[30][5] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19722_ (.D(_00052_),
    .Q(\CPU_Xreg_value_a4[30][6] ),
    .CLK(clknet_8_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19723_ (.D(_00053_),
    .Q(\CPU_Xreg_value_a4[30][7] ),
    .CLK(clknet_8_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19724_ (.D(_00054_),
    .Q(\CPU_Xreg_value_a4[30][8] ),
    .CLK(clknet_8_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19725_ (.D(_00055_),
    .Q(\CPU_Xreg_value_a4[30][9] ),
    .CLK(clknet_8_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19726_ (.D(_00056_),
    .Q(\CPU_Xreg_value_a4[30][10] ),
    .CLK(clknet_8_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19727_ (.D(_00057_),
    .Q(\CPU_Xreg_value_a4[30][11] ),
    .CLK(clknet_8_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19728_ (.D(_00058_),
    .Q(\CPU_Xreg_value_a4[30][12] ),
    .CLK(clknet_8_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19729_ (.D(_00059_),
    .Q(\CPU_Xreg_value_a4[30][13] ),
    .CLK(clknet_8_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19730_ (.D(_00060_),
    .Q(\CPU_Xreg_value_a4[30][14] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19731_ (.D(_00061_),
    .Q(\CPU_Xreg_value_a4[30][15] ),
    .CLK(clknet_8_36_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19732_ (.D(_00062_),
    .Q(\CPU_Xreg_value_a4[30][16] ),
    .CLK(clknet_8_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19733_ (.D(_00063_),
    .Q(\CPU_Xreg_value_a4[30][17] ),
    .CLK(clknet_8_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19734_ (.D(_00064_),
    .Q(\CPU_Xreg_value_a4[30][18] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19735_ (.D(_00065_),
    .Q(\CPU_Xreg_value_a4[30][19] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19736_ (.D(_00066_),
    .Q(\CPU_Xreg_value_a4[30][20] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19737_ (.D(_00067_),
    .Q(\CPU_Xreg_value_a4[30][21] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19738_ (.D(_00068_),
    .Q(\CPU_Xreg_value_a4[30][22] ),
    .CLK(clknet_8_176_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19739_ (.D(_00069_),
    .Q(\CPU_Xreg_value_a4[30][23] ),
    .CLK(clknet_8_176_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19740_ (.D(_00070_),
    .Q(\CPU_Xreg_value_a4[30][24] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19741_ (.D(_00071_),
    .Q(\CPU_Xreg_value_a4[30][25] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19742_ (.D(_00072_),
    .Q(\CPU_Xreg_value_a4[30][26] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19743_ (.D(_00073_),
    .Q(\CPU_Xreg_value_a4[30][27] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19744_ (.D(_00074_),
    .Q(\CPU_Xreg_value_a4[30][28] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19745_ (.D(_00075_),
    .Q(\CPU_Xreg_value_a4[30][29] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19746_ (.D(_00076_),
    .Q(\CPU_Xreg_value_a4[30][30] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19747_ (.D(_00077_),
    .Q(\CPU_Xreg_value_a4[30][31] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19748_ (.D(_00078_),
    .Q(\CPU_Xreg_value_a4[29][0] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19749_ (.D(_00079_),
    .Q(\CPU_Xreg_value_a4[29][1] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19750_ (.D(_00080_),
    .Q(\CPU_Xreg_value_a4[29][2] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19751_ (.D(_00081_),
    .Q(\CPU_Xreg_value_a4[29][3] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19752_ (.D(_00082_),
    .Q(\CPU_Xreg_value_a4[29][4] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19753_ (.D(_00083_),
    .Q(\CPU_Xreg_value_a4[29][5] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19754_ (.D(_00084_),
    .Q(\CPU_Xreg_value_a4[29][6] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19755_ (.D(_00085_),
    .Q(\CPU_Xreg_value_a4[29][7] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19756_ (.D(_00086_),
    .Q(\CPU_Xreg_value_a4[29][8] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19757_ (.D(_00087_),
    .Q(\CPU_Xreg_value_a4[29][9] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19758_ (.D(_00088_),
    .Q(\CPU_Xreg_value_a4[29][10] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19759_ (.D(_00089_),
    .Q(\CPU_Xreg_value_a4[29][11] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19760_ (.D(_00090_),
    .Q(\CPU_Xreg_value_a4[29][12] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19761_ (.D(_00091_),
    .Q(\CPU_Xreg_value_a4[29][13] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19762_ (.D(_00092_),
    .Q(\CPU_Xreg_value_a4[29][14] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19763_ (.D(_00093_),
    .Q(\CPU_Xreg_value_a4[29][15] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19764_ (.D(_00094_),
    .Q(\CPU_Xreg_value_a4[29][16] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19765_ (.D(_00095_),
    .Q(\CPU_Xreg_value_a4[29][17] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19766_ (.D(_00096_),
    .Q(\CPU_Xreg_value_a4[29][18] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19767_ (.D(_00097_),
    .Q(\CPU_Xreg_value_a4[29][19] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19768_ (.D(_00098_),
    .Q(\CPU_Xreg_value_a4[29][20] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19769_ (.D(_00099_),
    .Q(\CPU_Xreg_value_a4[29][21] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19770_ (.D(_00100_),
    .Q(\CPU_Xreg_value_a4[29][22] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19771_ (.D(_00101_),
    .Q(\CPU_Xreg_value_a4[29][23] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19772_ (.D(_00102_),
    .Q(\CPU_Xreg_value_a4[29][24] ),
    .CLK(clknet_8_163_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19773_ (.D(_00103_),
    .Q(\CPU_Xreg_value_a4[29][25] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19774_ (.D(_00104_),
    .Q(\CPU_Xreg_value_a4[29][26] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19775_ (.D(_00105_),
    .Q(\CPU_Xreg_value_a4[29][27] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19776_ (.D(_00106_),
    .Q(\CPU_Xreg_value_a4[29][28] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19777_ (.D(_00107_),
    .Q(\CPU_Xreg_value_a4[29][29] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19778_ (.D(_00108_),
    .Q(\CPU_Xreg_value_a4[29][30] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19779_ (.D(_00109_),
    .Q(\CPU_Xreg_value_a4[29][31] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19780_ (.D(_00110_),
    .Q(\CPU_Xreg_value_a4[28][0] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19781_ (.D(_00111_),
    .Q(\CPU_Xreg_value_a4[28][1] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19782_ (.D(_00112_),
    .Q(\CPU_Xreg_value_a4[28][2] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19783_ (.D(_00113_),
    .Q(\CPU_Xreg_value_a4[28][3] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19784_ (.D(_00114_),
    .Q(\CPU_Xreg_value_a4[28][4] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19785_ (.D(_00115_),
    .Q(\CPU_Xreg_value_a4[28][5] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19786_ (.D(_00116_),
    .Q(\CPU_Xreg_value_a4[28][6] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19787_ (.D(_00117_),
    .Q(\CPU_Xreg_value_a4[28][7] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19788_ (.D(_00118_),
    .Q(\CPU_Xreg_value_a4[28][8] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19789_ (.D(_00119_),
    .Q(\CPU_Xreg_value_a4[28][9] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19790_ (.D(_00120_),
    .Q(\CPU_Xreg_value_a4[28][10] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19791_ (.D(_00121_),
    .Q(\CPU_Xreg_value_a4[28][11] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19792_ (.D(_00122_),
    .Q(\CPU_Xreg_value_a4[28][12] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19793_ (.D(_00123_),
    .Q(\CPU_Xreg_value_a4[28][13] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19794_ (.D(_00124_),
    .Q(\CPU_Xreg_value_a4[28][14] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19795_ (.D(_00125_),
    .Q(\CPU_Xreg_value_a4[28][15] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19796_ (.D(_00126_),
    .Q(\CPU_Xreg_value_a4[28][16] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19797_ (.D(_00127_),
    .Q(\CPU_Xreg_value_a4[28][17] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19798_ (.D(_00128_),
    .Q(\CPU_Xreg_value_a4[28][18] ),
    .CLK(clknet_8_137_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19799_ (.D(_00129_),
    .Q(\CPU_Xreg_value_a4[28][19] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19800_ (.D(_00130_),
    .Q(\CPU_Xreg_value_a4[28][20] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19801_ (.D(_00131_),
    .Q(\CPU_Xreg_value_a4[28][21] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19802_ (.D(_00132_),
    .Q(\CPU_Xreg_value_a4[28][22] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19803_ (.D(_00133_),
    .Q(\CPU_Xreg_value_a4[28][23] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19804_ (.D(_00134_),
    .Q(\CPU_Xreg_value_a4[28][24] ),
    .CLK(clknet_8_163_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19805_ (.D(_00135_),
    .Q(\CPU_Xreg_value_a4[28][25] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19806_ (.D(_00136_),
    .Q(\CPU_Xreg_value_a4[28][26] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19807_ (.D(_00137_),
    .Q(\CPU_Xreg_value_a4[28][27] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19808_ (.D(_00138_),
    .Q(\CPU_Xreg_value_a4[28][28] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19809_ (.D(_00139_),
    .Q(\CPU_Xreg_value_a4[28][29] ),
    .CLK(clknet_8_166_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19810_ (.D(_00140_),
    .Q(\CPU_Xreg_value_a4[28][30] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19811_ (.D(_00141_),
    .Q(\CPU_Xreg_value_a4[28][31] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19812_ (.D(_00142_),
    .Q(\CPU_Xreg_value_a4[27][0] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19813_ (.D(_00143_),
    .Q(\CPU_Xreg_value_a4[27][1] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19814_ (.D(_00144_),
    .Q(\CPU_Xreg_value_a4[27][2] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19815_ (.D(_00145_),
    .Q(\CPU_Xreg_value_a4[27][3] ),
    .CLK(clknet_8_134_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19816_ (.D(_00146_),
    .Q(\CPU_Xreg_value_a4[27][4] ),
    .CLK(clknet_8_134_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19817_ (.D(_00147_),
    .Q(\CPU_Xreg_value_a4[27][5] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19818_ (.D(_00148_),
    .Q(\CPU_Xreg_value_a4[27][6] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19819_ (.D(_00149_),
    .Q(\CPU_Xreg_value_a4[27][7] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19820_ (.D(_00150_),
    .Q(\CPU_Xreg_value_a4[27][8] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19821_ (.D(_00151_),
    .Q(\CPU_Xreg_value_a4[27][9] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19822_ (.D(_00152_),
    .Q(\CPU_Xreg_value_a4[27][10] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19823_ (.D(_00153_),
    .Q(\CPU_Xreg_value_a4[27][11] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19824_ (.D(_00154_),
    .Q(\CPU_Xreg_value_a4[27][12] ),
    .CLK(clknet_8_9_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19825_ (.D(_00155_),
    .Q(\CPU_Xreg_value_a4[27][13] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19826_ (.D(_00156_),
    .Q(\CPU_Xreg_value_a4[27][14] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19827_ (.D(_00157_),
    .Q(\CPU_Xreg_value_a4[27][15] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19828_ (.D(_00158_),
    .Q(\CPU_Xreg_value_a4[27][16] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19829_ (.D(_00159_),
    .Q(\CPU_Xreg_value_a4[27][17] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19830_ (.D(_00160_),
    .Q(\CPU_Xreg_value_a4[27][18] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19831_ (.D(_00161_),
    .Q(\CPU_Xreg_value_a4[27][19] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19832_ (.D(_00162_),
    .Q(\CPU_Xreg_value_a4[27][20] ),
    .CLK(clknet_8_137_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19833_ (.D(_00163_),
    .Q(\CPU_Xreg_value_a4[27][21] ),
    .CLK(clknet_8_137_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19834_ (.D(_00164_),
    .Q(\CPU_Xreg_value_a4[27][22] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19835_ (.D(_00165_),
    .Q(\CPU_Xreg_value_a4[27][23] ),
    .CLK(clknet_8_161_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19836_ (.D(_00166_),
    .Q(\CPU_Xreg_value_a4[27][24] ),
    .CLK(clknet_8_163_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19837_ (.D(_00167_),
    .Q(\CPU_Xreg_value_a4[27][25] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19838_ (.D(_00168_),
    .Q(\CPU_Xreg_value_a4[27][26] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19839_ (.D(_00169_),
    .Q(\CPU_Xreg_value_a4[27][27] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19840_ (.D(_00170_),
    .Q(\CPU_Xreg_value_a4[27][28] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19841_ (.D(_00171_),
    .Q(\CPU_Xreg_value_a4[27][29] ),
    .CLK(clknet_8_169_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19842_ (.D(_00172_),
    .Q(\CPU_Xreg_value_a4[27][30] ),
    .CLK(clknet_8_137_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19843_ (.D(_00173_),
    .Q(\CPU_Xreg_value_a4[27][31] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19844_ (.D(_00174_),
    .Q(\CPU_Xreg_value_a4[26][0] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19845_ (.D(_00175_),
    .Q(\CPU_Xreg_value_a4[26][1] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19846_ (.D(_00176_),
    .Q(\CPU_Xreg_value_a4[26][2] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19847_ (.D(_00177_),
    .Q(\CPU_Xreg_value_a4[26][3] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19848_ (.D(_00178_),
    .Q(\CPU_Xreg_value_a4[26][4] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19849_ (.D(_00179_),
    .Q(\CPU_Xreg_value_a4[26][5] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19850_ (.D(_00180_),
    .Q(\CPU_Xreg_value_a4[26][6] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19851_ (.D(_00181_),
    .Q(\CPU_Xreg_value_a4[26][7] ),
    .CLK(clknet_8_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19852_ (.D(_00182_),
    .Q(\CPU_Xreg_value_a4[26][8] ),
    .CLK(clknet_8_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19853_ (.D(_00183_),
    .Q(\CPU_Xreg_value_a4[26][9] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19854_ (.D(_00184_),
    .Q(\CPU_Xreg_value_a4[26][10] ),
    .CLK(clknet_8_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19855_ (.D(_00185_),
    .Q(\CPU_Xreg_value_a4[26][11] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19856_ (.D(_00186_),
    .Q(\CPU_Xreg_value_a4[26][12] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19857_ (.D(_00187_),
    .Q(\CPU_Xreg_value_a4[26][13] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19858_ (.D(_00188_),
    .Q(\CPU_Xreg_value_a4[26][14] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19859_ (.D(_00189_),
    .Q(\CPU_Xreg_value_a4[26][15] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19860_ (.D(_00190_),
    .Q(\CPU_Xreg_value_a4[26][16] ),
    .CLK(clknet_8_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19861_ (.D(_00191_),
    .Q(\CPU_Xreg_value_a4[26][17] ),
    .CLK(clknet_8_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19862_ (.D(_00192_),
    .Q(\CPU_Xreg_value_a4[26][18] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19863_ (.D(_00193_),
    .Q(\CPU_Xreg_value_a4[26][19] ),
    .CLK(clknet_8_154_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19864_ (.D(_00194_),
    .Q(\CPU_Xreg_value_a4[26][20] ),
    .CLK(clknet_8_154_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19865_ (.D(_00195_),
    .Q(\CPU_Xreg_value_a4[26][21] ),
    .CLK(clknet_8_154_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19866_ (.D(_00196_),
    .Q(\CPU_Xreg_value_a4[26][22] ),
    .CLK(clknet_8_178_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19867_ (.D(_00197_),
    .Q(\CPU_Xreg_value_a4[26][23] ),
    .CLK(clknet_8_178_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19868_ (.D(_00198_),
    .Q(\CPU_Xreg_value_a4[26][24] ),
    .CLK(clknet_8_178_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19869_ (.D(_00199_),
    .Q(\CPU_Xreg_value_a4[26][25] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19870_ (.D(_00200_),
    .Q(\CPU_Xreg_value_a4[26][26] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19871_ (.D(_00201_),
    .Q(\CPU_Xreg_value_a4[26][27] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19872_ (.D(_00202_),
    .Q(\CPU_Xreg_value_a4[26][28] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19873_ (.D(_00203_),
    .Q(\CPU_Xreg_value_a4[26][29] ),
    .CLK(clknet_8_186_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19874_ (.D(_00204_),
    .Q(\CPU_Xreg_value_a4[26][30] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19875_ (.D(_00205_),
    .Q(\CPU_Xreg_value_a4[26][31] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19876_ (.D(_00206_),
    .Q(\CPU_Xreg_value_a4[25][0] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19877_ (.D(_00207_),
    .Q(\CPU_Xreg_value_a4[25][1] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19878_ (.D(_00208_),
    .Q(\CPU_Xreg_value_a4[25][2] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19879_ (.D(_00209_),
    .Q(\CPU_Xreg_value_a4[25][3] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19880_ (.D(_00210_),
    .Q(\CPU_Xreg_value_a4[25][4] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19881_ (.D(_00211_),
    .Q(\CPU_Xreg_value_a4[25][5] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19882_ (.D(_00212_),
    .Q(\CPU_Xreg_value_a4[25][6] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19883_ (.D(_00213_),
    .Q(\CPU_Xreg_value_a4[25][7] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19884_ (.D(_00214_),
    .Q(\CPU_Xreg_value_a4[25][8] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19885_ (.D(_00215_),
    .Q(\CPU_Xreg_value_a4[25][9] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19886_ (.D(_00216_),
    .Q(\CPU_Xreg_value_a4[25][10] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19887_ (.D(_00217_),
    .Q(\CPU_Xreg_value_a4[25][11] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19888_ (.D(_00218_),
    .Q(\CPU_Xreg_value_a4[25][12] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19889_ (.D(_00219_),
    .Q(\CPU_Xreg_value_a4[25][13] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19890_ (.D(_00220_),
    .Q(\CPU_Xreg_value_a4[25][14] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19891_ (.D(_00221_),
    .Q(\CPU_Xreg_value_a4[25][15] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19892_ (.D(_00222_),
    .Q(\CPU_Xreg_value_a4[25][16] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19893_ (.D(_00223_),
    .Q(\CPU_Xreg_value_a4[25][17] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19894_ (.D(_00224_),
    .Q(\CPU_Xreg_value_a4[25][18] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19895_ (.D(_00225_),
    .Q(\CPU_Xreg_value_a4[25][19] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19896_ (.D(_00226_),
    .Q(\CPU_Xreg_value_a4[25][20] ),
    .CLK(clknet_8_139_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19897_ (.D(_00227_),
    .Q(\CPU_Xreg_value_a4[25][21] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19898_ (.D(_00228_),
    .Q(\CPU_Xreg_value_a4[25][22] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19899_ (.D(_00229_),
    .Q(\CPU_Xreg_value_a4[25][23] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19900_ (.D(_00230_),
    .Q(\CPU_Xreg_value_a4[25][24] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19901_ (.D(_00231_),
    .Q(\CPU_Xreg_value_a4[25][25] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19902_ (.D(_00232_),
    .Q(\CPU_Xreg_value_a4[25][26] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19903_ (.D(_00233_),
    .Q(\CPU_Xreg_value_a4[25][27] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19904_ (.D(_00234_),
    .Q(\CPU_Xreg_value_a4[25][28] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19905_ (.D(_00235_),
    .Q(\CPU_Xreg_value_a4[25][29] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19906_ (.D(_00236_),
    .Q(\CPU_Xreg_value_a4[25][30] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19907_ (.D(_00237_),
    .Q(\CPU_Xreg_value_a4[25][31] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19908_ (.D(_00238_),
    .Q(\CPU_Xreg_value_a4[24][0] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19909_ (.D(_00239_),
    .Q(\CPU_Xreg_value_a4[24][1] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19910_ (.D(_00240_),
    .Q(\CPU_Xreg_value_a4[24][2] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19911_ (.D(_00241_),
    .Q(\CPU_Xreg_value_a4[24][3] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19912_ (.D(_00242_),
    .Q(\CPU_Xreg_value_a4[24][4] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19913_ (.D(_00243_),
    .Q(\CPU_Xreg_value_a4[24][5] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19914_ (.D(_00244_),
    .Q(\CPU_Xreg_value_a4[24][6] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19915_ (.D(_00245_),
    .Q(\CPU_Xreg_value_a4[24][7] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19916_ (.D(_00246_),
    .Q(\CPU_Xreg_value_a4[24][8] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19917_ (.D(_00247_),
    .Q(\CPU_Xreg_value_a4[24][9] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19918_ (.D(_00248_),
    .Q(\CPU_Xreg_value_a4[24][10] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19919_ (.D(_00249_),
    .Q(\CPU_Xreg_value_a4[24][11] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19920_ (.D(_00250_),
    .Q(\CPU_Xreg_value_a4[24][12] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19921_ (.D(_00251_),
    .Q(\CPU_Xreg_value_a4[24][13] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19922_ (.D(_00252_),
    .Q(\CPU_Xreg_value_a4[24][14] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19923_ (.D(_00253_),
    .Q(\CPU_Xreg_value_a4[24][15] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19924_ (.D(_00254_),
    .Q(\CPU_Xreg_value_a4[24][16] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19925_ (.D(_00255_),
    .Q(\CPU_Xreg_value_a4[24][17] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19926_ (.D(_00256_),
    .Q(\CPU_Xreg_value_a4[24][18] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19927_ (.D(_00257_),
    .Q(\CPU_Xreg_value_a4[24][19] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19928_ (.D(_00258_),
    .Q(\CPU_Xreg_value_a4[24][20] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19929_ (.D(_00259_),
    .Q(\CPU_Xreg_value_a4[24][21] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19930_ (.D(_00260_),
    .Q(\CPU_Xreg_value_a4[24][22] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19931_ (.D(_00261_),
    .Q(\CPU_Xreg_value_a4[24][23] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19932_ (.D(_00262_),
    .Q(\CPU_Xreg_value_a4[24][24] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19933_ (.D(_00263_),
    .Q(\CPU_Xreg_value_a4[24][25] ),
    .CLK(clknet_8_171_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19934_ (.D(_00264_),
    .Q(\CPU_Xreg_value_a4[24][26] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19935_ (.D(_00265_),
    .Q(\CPU_Xreg_value_a4[24][27] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19936_ (.D(_00266_),
    .Q(\CPU_Xreg_value_a4[24][28] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19937_ (.D(_00267_),
    .Q(\CPU_Xreg_value_a4[24][29] ),
    .CLK(clknet_8_163_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19938_ (.D(_00268_),
    .Q(\CPU_Xreg_value_a4[24][30] ),
    .CLK(clknet_8_163_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19939_ (.D(_00269_),
    .Q(\CPU_Xreg_value_a4[24][31] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19940_ (.D(_00270_),
    .Q(\CPU_Xreg_value_a4[23][0] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19941_ (.D(_00271_),
    .Q(\CPU_Xreg_value_a4[23][1] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19942_ (.D(_00272_),
    .Q(\CPU_Xreg_value_a4[23][2] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19943_ (.D(_00273_),
    .Q(\CPU_Xreg_value_a4[23][3] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19944_ (.D(_00274_),
    .Q(\CPU_Xreg_value_a4[23][4] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19945_ (.D(_00275_),
    .Q(\CPU_Xreg_value_a4[23][5] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19946_ (.D(_00276_),
    .Q(\CPU_Xreg_value_a4[23][6] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19947_ (.D(_00277_),
    .Q(\CPU_Xreg_value_a4[23][7] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19948_ (.D(_00278_),
    .Q(\CPU_Xreg_value_a4[23][8] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19949_ (.D(_00279_),
    .Q(\CPU_Xreg_value_a4[23][9] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19950_ (.D(_00280_),
    .Q(\CPU_Xreg_value_a4[23][10] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19951_ (.D(_00281_),
    .Q(\CPU_Xreg_value_a4[23][11] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19952_ (.D(_00282_),
    .Q(\CPU_Xreg_value_a4[23][12] ),
    .CLK(clknet_8_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19953_ (.D(_00283_),
    .Q(\CPU_Xreg_value_a4[23][13] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19954_ (.D(_00284_),
    .Q(\CPU_Xreg_value_a4[23][14] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19955_ (.D(_00285_),
    .Q(\CPU_Xreg_value_a4[23][15] ),
    .CLK(clknet_8_38_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19956_ (.D(_00286_),
    .Q(\CPU_Xreg_value_a4[23][16] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19957_ (.D(_00287_),
    .Q(\CPU_Xreg_value_a4[23][17] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19958_ (.D(_00288_),
    .Q(\CPU_Xreg_value_a4[23][18] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19959_ (.D(_00289_),
    .Q(\CPU_Xreg_value_a4[23][19] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19960_ (.D(_00290_),
    .Q(\CPU_Xreg_value_a4[23][20] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19961_ (.D(_00291_),
    .Q(\CPU_Xreg_value_a4[23][21] ),
    .CLK(clknet_8_143_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19962_ (.D(_00292_),
    .Q(\CPU_Xreg_value_a4[23][22] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19963_ (.D(_00293_),
    .Q(\CPU_Xreg_value_a4[23][23] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19964_ (.D(_00294_),
    .Q(\CPU_Xreg_value_a4[23][24] ),
    .CLK(clknet_8_167_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19965_ (.D(_00295_),
    .Q(\CPU_Xreg_value_a4[23][25] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19966_ (.D(_00296_),
    .Q(\CPU_Xreg_value_a4[23][26] ),
    .CLK(clknet_8_172_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19967_ (.D(_00297_),
    .Q(\CPU_Xreg_value_a4[23][27] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19968_ (.D(_00298_),
    .Q(\CPU_Xreg_value_a4[23][28] ),
    .CLK(clknet_8_172_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19969_ (.D(_00299_),
    .Q(\CPU_Xreg_value_a4[23][29] ),
    .CLK(clknet_8_172_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19970_ (.D(_00300_),
    .Q(\CPU_Xreg_value_a4[23][30] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19971_ (.D(_00301_),
    .Q(\CPU_Xreg_value_a4[23][31] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19972_ (.D(_00302_),
    .Q(\CPU_Xreg_value_a4[22][0] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19973_ (.D(_00303_),
    .Q(\CPU_Xreg_value_a4[22][1] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19974_ (.D(_00304_),
    .Q(\CPU_Xreg_value_a4[22][2] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19975_ (.D(_00305_),
    .Q(\CPU_Xreg_value_a4[22][3] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19976_ (.D(_00306_),
    .Q(\CPU_Xreg_value_a4[22][4] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19977_ (.D(_00307_),
    .Q(\CPU_Xreg_value_a4[22][5] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19978_ (.D(_00308_),
    .Q(\CPU_Xreg_value_a4[22][6] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19979_ (.D(_00309_),
    .Q(\CPU_Xreg_value_a4[22][7] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19980_ (.D(_00310_),
    .Q(\CPU_Xreg_value_a4[22][8] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19981_ (.D(_00311_),
    .Q(\CPU_Xreg_value_a4[22][9] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19982_ (.D(_00312_),
    .Q(\CPU_Xreg_value_a4[22][10] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19983_ (.D(_00313_),
    .Q(\CPU_Xreg_value_a4[22][11] ),
    .CLK(clknet_8_3_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19984_ (.D(_00314_),
    .Q(\CPU_Xreg_value_a4[22][12] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19985_ (.D(_00315_),
    .Q(\CPU_Xreg_value_a4[22][13] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19986_ (.D(_00316_),
    .Q(\CPU_Xreg_value_a4[22][14] ),
    .CLK(clknet_8_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19987_ (.D(_00317_),
    .Q(\CPU_Xreg_value_a4[22][15] ),
    .CLK(clknet_8_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19988_ (.D(_00318_),
    .Q(\CPU_Xreg_value_a4[22][16] ),
    .CLK(clknet_8_132_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19989_ (.D(_00319_),
    .Q(\CPU_Xreg_value_a4[22][17] ),
    .CLK(clknet_8_134_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19990_ (.D(_00320_),
    .Q(\CPU_Xreg_value_a4[22][18] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19991_ (.D(_00321_),
    .Q(\CPU_Xreg_value_a4[22][19] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19992_ (.D(_00322_),
    .Q(\CPU_Xreg_value_a4[22][20] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19993_ (.D(_00323_),
    .Q(\CPU_Xreg_value_a4[22][21] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19994_ (.D(_00324_),
    .Q(\CPU_Xreg_value_a4[22][22] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19995_ (.D(_00325_),
    .Q(\CPU_Xreg_value_a4[22][23] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19996_ (.D(_00326_),
    .Q(\CPU_Xreg_value_a4[22][24] ),
    .CLK(clknet_8_173_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19997_ (.D(_00327_),
    .Q(\CPU_Xreg_value_a4[22][25] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19998_ (.D(_00328_),
    .Q(\CPU_Xreg_value_a4[22][26] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _19999_ (.D(_00329_),
    .Q(\CPU_Xreg_value_a4[22][27] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20000_ (.D(_00330_),
    .Q(\CPU_Xreg_value_a4[22][28] ),
    .CLK(clknet_8_166_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20001_ (.D(_00331_),
    .Q(\CPU_Xreg_value_a4[22][29] ),
    .CLK(clknet_8_166_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20002_ (.D(_00332_),
    .Q(\CPU_Xreg_value_a4[22][30] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20003_ (.D(_00333_),
    .Q(\CPU_Xreg_value_a4[22][31] ),
    .CLK(clknet_8_134_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20004_ (.D(_00334_),
    .Q(\CPU_Xreg_value_a4[21][0] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20005_ (.D(_00335_),
    .Q(\CPU_Xreg_value_a4[21][1] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20006_ (.D(_00336_),
    .Q(\CPU_Xreg_value_a4[21][2] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20007_ (.D(_00337_),
    .Q(\CPU_Xreg_value_a4[21][3] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20008_ (.D(_00338_),
    .Q(\CPU_Xreg_value_a4[21][4] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20009_ (.D(_00339_),
    .Q(\CPU_Xreg_value_a4[21][5] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20010_ (.D(_00340_),
    .Q(\CPU_Xreg_value_a4[21][6] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20011_ (.D(_00341_),
    .Q(\CPU_Xreg_value_a4[21][7] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20012_ (.D(_00342_),
    .Q(\CPU_Xreg_value_a4[21][8] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20013_ (.D(_00343_),
    .Q(\CPU_Xreg_value_a4[21][9] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20014_ (.D(_00344_),
    .Q(\CPU_Xreg_value_a4[21][10] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20015_ (.D(_00345_),
    .Q(\CPU_Xreg_value_a4[21][11] ),
    .CLK(clknet_8_8_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20016_ (.D(_00346_),
    .Q(\CPU_Xreg_value_a4[21][12] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20017_ (.D(_00347_),
    .Q(\CPU_Xreg_value_a4[21][13] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20018_ (.D(_00348_),
    .Q(\CPU_Xreg_value_a4[21][14] ),
    .CLK(clknet_8_34_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20019_ (.D(_00349_),
    .Q(\CPU_Xreg_value_a4[21][15] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20020_ (.D(_00350_),
    .Q(\CPU_Xreg_value_a4[21][16] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20021_ (.D(_00351_),
    .Q(\CPU_Xreg_value_a4[21][17] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20022_ (.D(_00352_),
    .Q(\CPU_Xreg_value_a4[21][18] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20023_ (.D(_00353_),
    .Q(\CPU_Xreg_value_a4[21][19] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20024_ (.D(_00354_),
    .Q(\CPU_Xreg_value_a4[21][20] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20025_ (.D(_00355_),
    .Q(\CPU_Xreg_value_a4[21][21] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20026_ (.D(_00356_),
    .Q(\CPU_Xreg_value_a4[21][22] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20027_ (.D(_00357_),
    .Q(\CPU_Xreg_value_a4[21][23] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20028_ (.D(_00358_),
    .Q(\CPU_Xreg_value_a4[21][24] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20029_ (.D(_00359_),
    .Q(\CPU_Xreg_value_a4[21][25] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20030_ (.D(_00360_),
    .Q(\CPU_Xreg_value_a4[21][26] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20031_ (.D(_00361_),
    .Q(\CPU_Xreg_value_a4[21][27] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20032_ (.D(_00362_),
    .Q(\CPU_Xreg_value_a4[21][28] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20033_ (.D(_00363_),
    .Q(\CPU_Xreg_value_a4[21][29] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20034_ (.D(_00364_),
    .Q(\CPU_Xreg_value_a4[21][30] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20035_ (.D(_00365_),
    .Q(\CPU_Xreg_value_a4[21][31] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20036_ (.D(_00366_),
    .Q(\CPU_Xreg_value_a4[20][0] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20037_ (.D(_00367_),
    .Q(\CPU_Xreg_value_a4[20][1] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20038_ (.D(_00368_),
    .Q(\CPU_Xreg_value_a4[20][2] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20039_ (.D(_00369_),
    .Q(\CPU_Xreg_value_a4[20][3] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20040_ (.D(_00370_),
    .Q(\CPU_Xreg_value_a4[20][4] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20041_ (.D(_00371_),
    .Q(\CPU_Xreg_value_a4[20][5] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20042_ (.D(_00372_),
    .Q(\CPU_Xreg_value_a4[20][6] ),
    .CLK(clknet_8_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20043_ (.D(_00373_),
    .Q(\CPU_Xreg_value_a4[20][7] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20044_ (.D(_00374_),
    .Q(\CPU_Xreg_value_a4[20][8] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20045_ (.D(_00375_),
    .Q(\CPU_Xreg_value_a4[20][9] ),
    .CLK(clknet_8_0_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20046_ (.D(_00376_),
    .Q(\CPU_Xreg_value_a4[20][10] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20047_ (.D(_00377_),
    .Q(\CPU_Xreg_value_a4[20][11] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20048_ (.D(_00378_),
    .Q(\CPU_Xreg_value_a4[20][12] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20049_ (.D(_00379_),
    .Q(\CPU_Xreg_value_a4[20][13] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20050_ (.D(_00380_),
    .Q(\CPU_Xreg_value_a4[20][14] ),
    .CLK(clknet_8_32_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20051_ (.D(_00381_),
    .Q(\CPU_Xreg_value_a4[20][15] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20052_ (.D(_00382_),
    .Q(\CPU_Xreg_value_a4[20][16] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20053_ (.D(_00383_),
    .Q(\CPU_Xreg_value_a4[20][17] ),
    .CLK(clknet_8_130_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20054_ (.D(_00384_),
    .Q(\CPU_Xreg_value_a4[20][18] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20055_ (.D(_00385_),
    .Q(\CPU_Xreg_value_a4[20][19] ),
    .CLK(clknet_8_136_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20056_ (.D(_00386_),
    .Q(\CPU_Xreg_value_a4[20][20] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20057_ (.D(_00387_),
    .Q(\CPU_Xreg_value_a4[20][21] ),
    .CLK(clknet_8_138_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20058_ (.D(_00388_),
    .Q(\CPU_Xreg_value_a4[20][22] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20059_ (.D(_00389_),
    .Q(\CPU_Xreg_value_a4[20][23] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20060_ (.D(_00390_),
    .Q(\CPU_Xreg_value_a4[20][24] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20061_ (.D(_00391_),
    .Q(\CPU_Xreg_value_a4[20][25] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20062_ (.D(_00392_),
    .Q(\CPU_Xreg_value_a4[20][26] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20063_ (.D(_00393_),
    .Q(\CPU_Xreg_value_a4[20][27] ),
    .CLK(clknet_8_170_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20064_ (.D(_00394_),
    .Q(\CPU_Xreg_value_a4[20][28] ),
    .CLK(clknet_8_168_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20065_ (.D(_00395_),
    .Q(\CPU_Xreg_value_a4[20][29] ),
    .CLK(clknet_8_162_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20066_ (.D(_00396_),
    .Q(\CPU_Xreg_value_a4[20][30] ),
    .CLK(clknet_8_160_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20067_ (.D(_00397_),
    .Q(\CPU_Xreg_value_a4[20][31] ),
    .CLK(clknet_8_128_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20068_ (.D(_00398_),
    .Q(\CPU_Xreg_value_a4[19][0] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20069_ (.D(_00399_),
    .Q(\CPU_Xreg_value_a4[19][1] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20070_ (.D(_00400_),
    .Q(\CPU_Xreg_value_a4[19][2] ),
    .CLK(clknet_8_147_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20071_ (.D(_00401_),
    .Q(\CPU_Xreg_value_a4[19][3] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20072_ (.D(_00402_),
    .Q(\CPU_Xreg_value_a4[19][4] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20073_ (.D(_00403_),
    .Q(\CPU_Xreg_value_a4[19][5] ),
    .CLK(clknet_8_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20074_ (.D(_00404_),
    .Q(\CPU_Xreg_value_a4[19][6] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20075_ (.D(_00405_),
    .Q(\CPU_Xreg_value_a4[19][7] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20076_ (.D(_00406_),
    .Q(\CPU_Xreg_value_a4[19][8] ),
    .CLK(clknet_8_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20077_ (.D(_00407_),
    .Q(\CPU_Xreg_value_a4[19][9] ),
    .CLK(clknet_8_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20078_ (.D(_00408_),
    .Q(\CPU_Xreg_value_a4[19][10] ),
    .CLK(clknet_8_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20079_ (.D(_00409_),
    .Q(\CPU_Xreg_value_a4[19][11] ),
    .CLK(clknet_8_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20080_ (.D(_00410_),
    .Q(\CPU_Xreg_value_a4[19][12] ),
    .CLK(clknet_8_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20081_ (.D(_00411_),
    .Q(\CPU_Xreg_value_a4[19][13] ),
    .CLK(clknet_8_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20082_ (.D(_00412_),
    .Q(\CPU_Xreg_value_a4[19][14] ),
    .CLK(clknet_8_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20083_ (.D(_00413_),
    .Q(\CPU_Xreg_value_a4[19][15] ),
    .CLK(clknet_8_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20084_ (.D(_00414_),
    .Q(\CPU_Xreg_value_a4[19][16] ),
    .CLK(clknet_8_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20085_ (.D(_00415_),
    .Q(\CPU_Xreg_value_a4[19][17] ),
    .CLK(clknet_8_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20086_ (.D(_00416_),
    .Q(\CPU_Xreg_value_a4[19][18] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20087_ (.D(_00417_),
    .Q(\CPU_Xreg_value_a4[19][19] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20088_ (.D(_00418_),
    .Q(\CPU_Xreg_value_a4[19][20] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20089_ (.D(_00419_),
    .Q(\CPU_Xreg_value_a4[19][21] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20090_ (.D(_00420_),
    .Q(\CPU_Xreg_value_a4[19][22] ),
    .CLK(clknet_8_177_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20091_ (.D(_00421_),
    .Q(\CPU_Xreg_value_a4[19][23] ),
    .CLK(clknet_8_177_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20092_ (.D(_00422_),
    .Q(\CPU_Xreg_value_a4[19][24] ),
    .CLK(clknet_8_182_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20093_ (.D(_00423_),
    .Q(\CPU_Xreg_value_a4[19][25] ),
    .CLK(clknet_8_182_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20094_ (.D(_00424_),
    .Q(\CPU_Xreg_value_a4[19][26] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20095_ (.D(_00425_),
    .Q(\CPU_Xreg_value_a4[19][27] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20096_ (.D(_00426_),
    .Q(\CPU_Xreg_value_a4[19][28] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20097_ (.D(_00427_),
    .Q(\CPU_Xreg_value_a4[19][29] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20098_ (.D(_00428_),
    .Q(\CPU_Xreg_value_a4[19][30] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20099_ (.D(_00429_),
    .Q(\CPU_Xreg_value_a4[19][31] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20100_ (.D(_00430_),
    .Q(\CPU_Xreg_value_a4[18][0] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20101_ (.D(_00431_),
    .Q(\CPU_Xreg_value_a4[18][1] ),
    .CLK(clknet_8_42_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20102_ (.D(_00432_),
    .Q(\CPU_Xreg_value_a4[18][2] ),
    .CLK(clknet_8_129_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20103_ (.D(_00433_),
    .Q(\CPU_Xreg_value_a4[18][3] ),
    .CLK(clknet_8_40_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20104_ (.D(_00434_),
    .Q(\CPU_Xreg_value_a4[18][4] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20105_ (.D(_00435_),
    .Q(\CPU_Xreg_value_a4[18][5] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20106_ (.D(_00436_),
    .Q(\CPU_Xreg_value_a4[18][6] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20107_ (.D(_00437_),
    .Q(\CPU_Xreg_value_a4[18][7] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20108_ (.D(_00438_),
    .Q(\CPU_Xreg_value_a4[18][8] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20109_ (.D(_00439_),
    .Q(\CPU_Xreg_value_a4[18][9] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20110_ (.D(_00440_),
    .Q(\CPU_Xreg_value_a4[18][10] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20111_ (.D(_00441_),
    .Q(\CPU_Xreg_value_a4[18][11] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20112_ (.D(_00442_),
    .Q(\CPU_Xreg_value_a4[18][12] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20113_ (.D(_00443_),
    .Q(\CPU_Xreg_value_a4[18][13] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20114_ (.D(_00444_),
    .Q(\CPU_Xreg_value_a4[18][14] ),
    .CLK(clknet_8_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20115_ (.D(_00445_),
    .Q(\CPU_Xreg_value_a4[18][15] ),
    .CLK(clknet_8_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20116_ (.D(_00446_),
    .Q(\CPU_Xreg_value_a4[18][16] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20117_ (.D(_00447_),
    .Q(\CPU_Xreg_value_a4[18][17] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20118_ (.D(_00448_),
    .Q(\CPU_Xreg_value_a4[18][18] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20119_ (.D(_00449_),
    .Q(\CPU_Xreg_value_a4[18][19] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20120_ (.D(_00450_),
    .Q(\CPU_Xreg_value_a4[18][20] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20121_ (.D(_00451_),
    .Q(\CPU_Xreg_value_a4[18][21] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20122_ (.D(_00452_),
    .Q(\CPU_Xreg_value_a4[18][22] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20123_ (.D(_00453_),
    .Q(\CPU_Xreg_value_a4[18][23] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20124_ (.D(_00454_),
    .Q(\CPU_Xreg_value_a4[18][24] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20125_ (.D(_00455_),
    .Q(\CPU_Xreg_value_a4[18][25] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20126_ (.D(_00456_),
    .Q(\CPU_Xreg_value_a4[18][26] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20127_ (.D(_00457_),
    .Q(\CPU_Xreg_value_a4[18][27] ),
    .CLK(clknet_8_174_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20128_ (.D(_00458_),
    .Q(\CPU_Xreg_value_a4[18][28] ),
    .CLK(clknet_8_172_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20129_ (.D(_00459_),
    .Q(\CPU_Xreg_value_a4[18][29] ),
    .CLK(clknet_8_172_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20130_ (.D(_00460_),
    .Q(\CPU_Xreg_value_a4[18][30] ),
    .CLK(clknet_8_137_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20131_ (.D(_00461_),
    .Q(\CPU_Xreg_value_a4[18][31] ),
    .CLK(clknet_8_131_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20132_ (.D(_00462_),
    .Q(\CPU_Xreg_value_a4[17][0] ),
    .CLK(clknet_8_133_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20133_ (.D(_00463_),
    .Q(\CPU_Xreg_value_a4[17][1] ),
    .CLK(clknet_8_43_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20134_ (.D(_00464_),
    .Q(\CPU_Xreg_value_a4[17][2] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20135_ (.D(_00465_),
    .Q(\CPU_Xreg_value_a4[17][3] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20136_ (.D(_00466_),
    .Q(\CPU_Xreg_value_a4[17][4] ),
    .CLK(clknet_8_46_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20137_ (.D(_00467_),
    .Q(\CPU_Xreg_value_a4[17][5] ),
    .CLK(clknet_8_44_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20138_ (.D(_00468_),
    .Q(\CPU_Xreg_value_a4[17][6] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20139_ (.D(_00469_),
    .Q(\CPU_Xreg_value_a4[17][7] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20140_ (.D(_00470_),
    .Q(\CPU_Xreg_value_a4[17][8] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20141_ (.D(_00471_),
    .Q(\CPU_Xreg_value_a4[17][9] ),
    .CLK(clknet_8_1_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20142_ (.D(_00472_),
    .Q(\CPU_Xreg_value_a4[17][10] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20143_ (.D(_00473_),
    .Q(\CPU_Xreg_value_a4[17][11] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20144_ (.D(_00474_),
    .Q(\CPU_Xreg_value_a4[17][12] ),
    .CLK(clknet_8_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20145_ (.D(_00475_),
    .Q(\CPU_Xreg_value_a4[17][13] ),
    .CLK(clknet_8_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20146_ (.D(_00476_),
    .Q(\CPU_Xreg_value_a4[17][14] ),
    .CLK(clknet_8_33_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20147_ (.D(_00477_),
    .Q(\CPU_Xreg_value_a4[17][15] ),
    .CLK(clknet_8_35_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20148_ (.D(_00478_),
    .Q(\CPU_Xreg_value_a4[17][16] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20149_ (.D(_00479_),
    .Q(\CPU_Xreg_value_a4[17][17] ),
    .CLK(clknet_8_41_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20150_ (.D(_00480_),
    .Q(\CPU_Xreg_value_a4[17][18] ),
    .CLK(clknet_8_141_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20151_ (.D(_00481_),
    .Q(\CPU_Xreg_value_a4[17][19] ),
    .CLK(clknet_8_140_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20152_ (.D(_00482_),
    .Q(\CPU_Xreg_value_a4[17][20] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20153_ (.D(_00483_),
    .Q(\CPU_Xreg_value_a4[17][21] ),
    .CLK(clknet_8_142_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20154_ (.D(_00484_),
    .Q(\CPU_Xreg_value_a4[17][22] ),
    .CLK(clknet_8_165_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20155_ (.D(_00485_),
    .Q(\CPU_Xreg_value_a4[17][23] ),
    .CLK(clknet_8_164_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20156_ (.D(_00486_),
    .Q(\CPU_Xreg_value_a4[17][24] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20157_ (.D(_00487_),
    .Q(\CPU_Xreg_value_a4[17][25] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20158_ (.D(_00488_),
    .Q(\CPU_Xreg_value_a4[17][26] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20159_ (.D(_00489_),
    .Q(\CPU_Xreg_value_a4[17][27] ),
    .CLK(clknet_8_175_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20160_ (.D(_00490_),
    .Q(\CPU_Xreg_value_a4[17][28] ),
    .CLK(clknet_8_166_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20161_ (.D(_00491_),
    .Q(\CPU_Xreg_value_a4[17][29] ),
    .CLK(clknet_8_166_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20162_ (.D(_00492_),
    .Q(\CPU_Xreg_value_a4[17][30] ),
    .CLK(clknet_8_135_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20163_ (.D(_00493_),
    .Q(\CPU_Xreg_value_a4[17][31] ),
    .CLK(clknet_8_134_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20164_ (.D(_00494_),
    .Q(\CPU_Xreg_value_a4[16][0] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20165_ (.D(_00495_),
    .Q(\CPU_Xreg_value_a4[16][1] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20166_ (.D(_00496_),
    .Q(\CPU_Xreg_value_a4[16][2] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20167_ (.D(_00497_),
    .Q(\CPU_Xreg_value_a4[16][3] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20168_ (.D(_00498_),
    .Q(\CPU_Xreg_value_a4[16][4] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20169_ (.D(_00499_),
    .Q(\CPU_Xreg_value_a4[16][5] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20170_ (.D(_00500_),
    .Q(\CPU_Xreg_value_a4[16][6] ),
    .CLK(clknet_8_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20171_ (.D(_00501_),
    .Q(\CPU_Xreg_value_a4[16][7] ),
    .CLK(clknet_8_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20172_ (.D(_00502_),
    .Q(\CPU_Xreg_value_a4[16][8] ),
    .CLK(clknet_8_12_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20173_ (.D(_00503_),
    .Q(\CPU_Xreg_value_a4[16][9] ),
    .CLK(clknet_8_14_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20174_ (.D(_00504_),
    .Q(\CPU_Xreg_value_a4[16][10] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20175_ (.D(_00505_),
    .Q(\CPU_Xreg_value_a4[16][11] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20176_ (.D(_00506_),
    .Q(\CPU_Xreg_value_a4[16][12] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20177_ (.D(_00507_),
    .Q(\CPU_Xreg_value_a4[16][13] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20178_ (.D(_00508_),
    .Q(\CPU_Xreg_value_a4[16][14] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20179_ (.D(_00509_),
    .Q(\CPU_Xreg_value_a4[16][15] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20180_ (.D(_00510_),
    .Q(\CPU_Xreg_value_a4[16][16] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20181_ (.D(_00511_),
    .Q(\CPU_Xreg_value_a4[16][17] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20182_ (.D(_00512_),
    .Q(\CPU_Xreg_value_a4[16][18] ),
    .CLK(clknet_8_152_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20183_ (.D(_00513_),
    .Q(\CPU_Xreg_value_a4[16][19] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20184_ (.D(_00514_),
    .Q(\CPU_Xreg_value_a4[16][20] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20185_ (.D(_00515_),
    .Q(\CPU_Xreg_value_a4[16][21] ),
    .CLK(clknet_8_153_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20186_ (.D(_00516_),
    .Q(\CPU_Xreg_value_a4[16][22] ),
    .CLK(clknet_8_176_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20187_ (.D(_00517_),
    .Q(\CPU_Xreg_value_a4[16][23] ),
    .CLK(clknet_8_178_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20188_ (.D(_00518_),
    .Q(\CPU_Xreg_value_a4[16][24] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20189_ (.D(_00519_),
    .Q(\CPU_Xreg_value_a4[16][25] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20190_ (.D(_00520_),
    .Q(\CPU_Xreg_value_a4[16][26] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20191_ (.D(_00521_),
    .Q(\CPU_Xreg_value_a4[16][27] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20192_ (.D(_00522_),
    .Q(\CPU_Xreg_value_a4[16][28] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20193_ (.D(_00523_),
    .Q(\CPU_Xreg_value_a4[16][29] ),
    .CLK(clknet_8_184_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20194_ (.D(_00524_),
    .Q(\CPU_Xreg_value_a4[16][30] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20195_ (.D(_00525_),
    .Q(\CPU_Xreg_value_a4[16][31] ),
    .CLK(clknet_8_146_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20196_ (.D(_00526_),
    .Q(\CPU_Xreg_value_a4[15][0] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20197_ (.D(_00527_),
    .Q(\CPU_Xreg_value_a4[15][1] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20198_ (.D(_00528_),
    .Q(\CPU_Xreg_value_a4[15][2] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20199_ (.D(_00529_),
    .Q(\CPU_Xreg_value_a4[15][3] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20200_ (.D(_00530_),
    .Q(\CPU_Xreg_value_a4[15][4] ),
    .CLK(clknet_8_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20201_ (.D(_00531_),
    .Q(\CPU_Xreg_value_a4[15][5] ),
    .CLK(clknet_8_57_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20202_ (.D(_00532_),
    .Q(\CPU_Xreg_value_a4[15][6] ),
    .CLK(clknet_8_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20203_ (.D(_00533_),
    .Q(\CPU_Xreg_value_a4[15][7] ),
    .CLK(clknet_8_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20204_ (.D(_00534_),
    .Q(\CPU_Xreg_value_a4[15][8] ),
    .CLK(clknet_8_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20205_ (.D(_00535_),
    .Q(\CPU_Xreg_value_a4[15][9] ),
    .CLK(clknet_8_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20206_ (.D(_00536_),
    .Q(\CPU_Xreg_value_a4[15][10] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20207_ (.D(_00537_),
    .Q(\CPU_Xreg_value_a4[15][11] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20208_ (.D(_00538_),
    .Q(\CPU_Xreg_value_a4[15][12] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20209_ (.D(_00539_),
    .Q(\CPU_Xreg_value_a4[15][13] ),
    .CLK(clknet_8_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20210_ (.D(_00540_),
    .Q(\CPU_Xreg_value_a4[15][14] ),
    .CLK(clknet_8_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20211_ (.D(_00541_),
    .Q(\CPU_Xreg_value_a4[15][15] ),
    .CLK(clknet_8_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20212_ (.D(_00542_),
    .Q(\CPU_Xreg_value_a4[15][16] ),
    .CLK(clknet_8_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20213_ (.D(_00543_),
    .Q(\CPU_Xreg_value_a4[15][17] ),
    .CLK(clknet_8_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20214_ (.D(_00544_),
    .Q(\CPU_Xreg_value_a4[15][18] ),
    .CLK(clknet_8_156_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20215_ (.D(_00545_),
    .Q(\CPU_Xreg_value_a4[15][19] ),
    .CLK(clknet_8_156_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20216_ (.D(_00546_),
    .Q(\CPU_Xreg_value_a4[15][20] ),
    .CLK(clknet_8_156_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20217_ (.D(_00547_),
    .Q(\CPU_Xreg_value_a4[15][21] ),
    .CLK(clknet_8_156_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20218_ (.D(_00548_),
    .Q(\CPU_Xreg_value_a4[15][22] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20219_ (.D(_00549_),
    .Q(\CPU_Xreg_value_a4[15][23] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20220_ (.D(_00550_),
    .Q(\CPU_Xreg_value_a4[15][24] ),
    .CLK(clknet_8_182_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20221_ (.D(_00551_),
    .Q(\CPU_Xreg_value_a4[15][25] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20222_ (.D(_00552_),
    .Q(\CPU_Xreg_value_a4[15][26] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20223_ (.D(_00553_),
    .Q(\CPU_Xreg_value_a4[15][27] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20224_ (.D(_00554_),
    .Q(\CPU_Xreg_value_a4[15][28] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20225_ (.D(_00555_),
    .Q(\CPU_Xreg_value_a4[15][29] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20226_ (.D(_00556_),
    .Q(\CPU_Xreg_value_a4[15][30] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20227_ (.D(_00557_),
    .Q(\CPU_Xreg_value_a4[15][31] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20228_ (.D(_00558_),
    .Q(\CPU_Xreg_value_a4[14][0] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20229_ (.D(_00559_),
    .Q(\CPU_Xreg_value_a4[14][1] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20230_ (.D(_00560_),
    .Q(\CPU_Xreg_value_a4[14][2] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20231_ (.D(_00561_),
    .Q(\CPU_Xreg_value_a4[14][3] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20232_ (.D(_00562_),
    .Q(\CPU_Xreg_value_a4[14][4] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20233_ (.D(_00563_),
    .Q(\CPU_Xreg_value_a4[14][5] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20234_ (.D(_00564_),
    .Q(\CPU_Xreg_value_a4[14][6] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20235_ (.D(_00565_),
    .Q(\CPU_Xreg_value_a4[14][7] ),
    .CLK(clknet_8_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20236_ (.D(_00566_),
    .Q(\CPU_Xreg_value_a4[14][8] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20237_ (.D(_00567_),
    .Q(\CPU_Xreg_value_a4[14][9] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20238_ (.D(_00568_),
    .Q(\CPU_Xreg_value_a4[14][10] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20239_ (.D(_00569_),
    .Q(\CPU_Xreg_value_a4[14][11] ),
    .CLK(clknet_8_4_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20240_ (.D(_00570_),
    .Q(\CPU_Xreg_value_a4[14][12] ),
    .CLK(clknet_8_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20241_ (.D(_00571_),
    .Q(\CPU_Xreg_value_a4[14][13] ),
    .CLK(clknet_8_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20242_ (.D(_00572_),
    .Q(\CPU_Xreg_value_a4[14][14] ),
    .CLK(clknet_8_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20243_ (.D(_00573_),
    .Q(\CPU_Xreg_value_a4[14][15] ),
    .CLK(clknet_8_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20244_ (.D(_00574_),
    .Q(\CPU_Xreg_value_a4[14][16] ),
    .CLK(clknet_8_51_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20245_ (.D(_00575_),
    .Q(\CPU_Xreg_value_a4[14][17] ),
    .CLK(clknet_8_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20246_ (.D(_00576_),
    .Q(\CPU_Xreg_value_a4[14][18] ),
    .CLK(clknet_8_156_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20247_ (.D(_00577_),
    .Q(\CPU_Xreg_value_a4[14][19] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20248_ (.D(_00578_),
    .Q(\CPU_Xreg_value_a4[14][20] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20249_ (.D(_00579_),
    .Q(\CPU_Xreg_value_a4[14][21] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20250_ (.D(_00580_),
    .Q(\CPU_Xreg_value_a4[14][22] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20251_ (.D(_00581_),
    .Q(\CPU_Xreg_value_a4[14][23] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20252_ (.D(_00582_),
    .Q(\CPU_Xreg_value_a4[14][24] ),
    .CLK(clknet_8_182_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20253_ (.D(_00583_),
    .Q(\CPU_Xreg_value_a4[14][25] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20254_ (.D(_00584_),
    .Q(\CPU_Xreg_value_a4[14][26] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20255_ (.D(_00585_),
    .Q(\CPU_Xreg_value_a4[14][27] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20256_ (.D(_00586_),
    .Q(\CPU_Xreg_value_a4[14][28] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20257_ (.D(_00587_),
    .Q(\CPU_Xreg_value_a4[14][29] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20258_ (.D(_00588_),
    .Q(\CPU_Xreg_value_a4[14][30] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20259_ (.D(_00589_),
    .Q(\CPU_Xreg_value_a4[14][31] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20260_ (.D(_00590_),
    .Q(\CPU_Xreg_value_a4[13][0] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20261_ (.D(_00591_),
    .Q(\CPU_Xreg_value_a4[13][1] ),
    .CLK(clknet_8_47_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20262_ (.D(_00592_),
    .Q(\CPU_Xreg_value_a4[13][2] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20263_ (.D(_00593_),
    .Q(\CPU_Xreg_value_a4[13][3] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20264_ (.D(_00594_),
    .Q(\CPU_Xreg_value_a4[13][4] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20265_ (.D(_00595_),
    .Q(\CPU_Xreg_value_a4[13][5] ),
    .CLK(clknet_8_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20266_ (.D(_00596_),
    .Q(\CPU_Xreg_value_a4[13][6] ),
    .CLK(clknet_8_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20267_ (.D(_00597_),
    .Q(\CPU_Xreg_value_a4[13][7] ),
    .CLK(clknet_8_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20268_ (.D(_00598_),
    .Q(\CPU_Xreg_value_a4[13][8] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20269_ (.D(_00599_),
    .Q(\CPU_Xreg_value_a4[13][9] ),
    .CLK(clknet_8_6_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20270_ (.D(_00600_),
    .Q(\CPU_Xreg_value_a4[13][10] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20271_ (.D(_00601_),
    .Q(\CPU_Xreg_value_a4[13][11] ),
    .CLK(clknet_8_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20272_ (.D(_00602_),
    .Q(\CPU_Xreg_value_a4[13][12] ),
    .CLK(clknet_8_13_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20273_ (.D(_00603_),
    .Q(\CPU_Xreg_value_a4[13][13] ),
    .CLK(clknet_8_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20274_ (.D(_00604_),
    .Q(\CPU_Xreg_value_a4[13][14] ),
    .CLK(clknet_8_54_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20275_ (.D(_00605_),
    .Q(\CPU_Xreg_value_a4[13][15] ),
    .CLK(clknet_8_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20276_ (.D(_00606_),
    .Q(\CPU_Xreg_value_a4[13][16] ),
    .CLK(clknet_8_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20277_ (.D(_00607_),
    .Q(\CPU_Xreg_value_a4[13][17] ),
    .CLK(clknet_8_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20278_ (.D(_00608_),
    .Q(\CPU_Xreg_value_a4[13][18] ),
    .CLK(clknet_8_45_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20279_ (.D(_00609_),
    .Q(\CPU_Xreg_value_a4[13][19] ),
    .CLK(clknet_8_154_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20280_ (.D(_00610_),
    .Q(\CPU_Xreg_value_a4[13][20] ),
    .CLK(clknet_8_155_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20281_ (.D(_00611_),
    .Q(\CPU_Xreg_value_a4[13][21] ),
    .CLK(clknet_8_155_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20282_ (.D(_00612_),
    .Q(\CPU_Xreg_value_a4[13][22] ),
    .CLK(clknet_8_176_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20283_ (.D(_00613_),
    .Q(\CPU_Xreg_value_a4[13][23] ),
    .CLK(clknet_8_176_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20284_ (.D(_00614_),
    .Q(\CPU_Xreg_value_a4[13][24] ),
    .CLK(clknet_8_179_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20285_ (.D(_00615_),
    .Q(\CPU_Xreg_value_a4[13][25] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20286_ (.D(_00616_),
    .Q(\CPU_Xreg_value_a4[13][26] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20287_ (.D(_00617_),
    .Q(\CPU_Xreg_value_a4[13][27] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20288_ (.D(_00618_),
    .Q(\CPU_Xreg_value_a4[13][28] ),
    .CLK(clknet_8_185_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20289_ (.D(_00619_),
    .Q(\CPU_Xreg_value_a4[13][29] ),
    .CLK(clknet_8_185_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20290_ (.D(_00620_),
    .Q(\CPU_Xreg_value_a4[13][30] ),
    .CLK(clknet_8_179_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20291_ (.D(_00621_),
    .Q(\CPU_Xreg_value_a4[13][31] ),
    .CLK(clknet_8_147_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20292_ (.D(_00622_),
    .Q(\CPU_Xreg_value_a4[12][0] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20293_ (.D(_00623_),
    .Q(\CPU_Xreg_value_a4[12][1] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20294_ (.D(_00624_),
    .Q(\CPU_Xreg_value_a4[12][2] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20295_ (.D(_00625_),
    .Q(\CPU_Xreg_value_a4[12][3] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20296_ (.D(_00626_),
    .Q(\CPU_Xreg_value_a4[12][4] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20297_ (.D(_00627_),
    .Q(\CPU_Xreg_value_a4[12][5] ),
    .CLK(clknet_8_59_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20298_ (.D(_00628_),
    .Q(\CPU_Xreg_value_a4[12][6] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20299_ (.D(_00629_),
    .Q(\CPU_Xreg_value_a4[12][7] ),
    .CLK(clknet_8_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20300_ (.D(_00630_),
    .Q(\CPU_Xreg_value_a4[12][8] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20301_ (.D(_00631_),
    .Q(\CPU_Xreg_value_a4[12][9] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20302_ (.D(_00632_),
    .Q(\CPU_Xreg_value_a4[12][10] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20303_ (.D(_00633_),
    .Q(\CPU_Xreg_value_a4[12][11] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20304_ (.D(_00634_),
    .Q(\CPU_Xreg_value_a4[12][12] ),
    .CLK(clknet_8_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20305_ (.D(_00635_),
    .Q(\CPU_Xreg_value_a4[12][13] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20306_ (.D(_00636_),
    .Q(\CPU_Xreg_value_a4[12][14] ),
    .CLK(clknet_8_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20307_ (.D(_00637_),
    .Q(\CPU_Xreg_value_a4[12][15] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20308_ (.D(_00638_),
    .Q(\CPU_Xreg_value_a4[12][16] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20309_ (.D(_00639_),
    .Q(\CPU_Xreg_value_a4[12][17] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20310_ (.D(_00640_),
    .Q(\CPU_Xreg_value_a4[12][18] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20311_ (.D(_00641_),
    .Q(\CPU_Xreg_value_a4[12][19] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20312_ (.D(_00642_),
    .Q(\CPU_Xreg_value_a4[12][20] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20313_ (.D(_00643_),
    .Q(\CPU_Xreg_value_a4[12][21] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20314_ (.D(_00644_),
    .Q(\CPU_Xreg_value_a4[12][22] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20315_ (.D(_00645_),
    .Q(\CPU_Xreg_value_a4[12][23] ),
    .CLK(clknet_8_183_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20316_ (.D(_00646_),
    .Q(\CPU_Xreg_value_a4[12][24] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20317_ (.D(_00647_),
    .Q(\CPU_Xreg_value_a4[12][25] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20318_ (.D(_00648_),
    .Q(\CPU_Xreg_value_a4[12][26] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20319_ (.D(_00649_),
    .Q(\CPU_Xreg_value_a4[12][27] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20320_ (.D(_00650_),
    .Q(\CPU_Xreg_value_a4[12][28] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20321_ (.D(_00651_),
    .Q(\CPU_Xreg_value_a4[12][29] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20322_ (.D(_00652_),
    .Q(\CPU_Xreg_value_a4[12][30] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20323_ (.D(_00653_),
    .Q(\CPU_Xreg_value_a4[12][31] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20324_ (.D(_00654_),
    .Q(\CPU_Xreg_value_a4[11][0] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20325_ (.D(_00655_),
    .Q(\CPU_Xreg_value_a4[11][1] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20326_ (.D(_00656_),
    .Q(\CPU_Xreg_value_a4[11][2] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20327_ (.D(_00657_),
    .Q(\CPU_Xreg_value_a4[11][3] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20328_ (.D(_00658_),
    .Q(\CPU_Xreg_value_a4[11][4] ),
    .CLK(clknet_8_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20329_ (.D(_00659_),
    .Q(\CPU_Xreg_value_a4[11][5] ),
    .CLK(clknet_8_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20330_ (.D(_00660_),
    .Q(\CPU_Xreg_value_a4[11][6] ),
    .CLK(clknet_8_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20331_ (.D(_00661_),
    .Q(\CPU_Xreg_value_a4[11][7] ),
    .CLK(clknet_8_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20332_ (.D(_00662_),
    .Q(\CPU_Xreg_value_a4[11][8] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20333_ (.D(_00663_),
    .Q(\CPU_Xreg_value_a4[11][9] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20334_ (.D(_00664_),
    .Q(\CPU_Xreg_value_a4[11][10] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20335_ (.D(_00665_),
    .Q(\CPU_Xreg_value_a4[11][11] ),
    .CLK(clknet_8_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20336_ (.D(_00666_),
    .Q(\CPU_Xreg_value_a4[11][12] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20337_ (.D(_00667_),
    .Q(\CPU_Xreg_value_a4[11][13] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20338_ (.D(_00668_),
    .Q(\CPU_Xreg_value_a4[11][14] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20339_ (.D(_00669_),
    .Q(\CPU_Xreg_value_a4[11][15] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20340_ (.D(_00670_),
    .Q(\CPU_Xreg_value_a4[11][16] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20341_ (.D(_00671_),
    .Q(\CPU_Xreg_value_a4[11][17] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20342_ (.D(_00672_),
    .Q(\CPU_Xreg_value_a4[11][18] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20343_ (.D(_00673_),
    .Q(\CPU_Xreg_value_a4[11][19] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20344_ (.D(_00674_),
    .Q(\CPU_Xreg_value_a4[11][20] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20345_ (.D(_00675_),
    .Q(\CPU_Xreg_value_a4[11][21] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20346_ (.D(_00676_),
    .Q(\CPU_Xreg_value_a4[11][22] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20347_ (.D(_00677_),
    .Q(\CPU_Xreg_value_a4[11][23] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20348_ (.D(_00678_),
    .Q(\CPU_Xreg_value_a4[11][24] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20349_ (.D(_00679_),
    .Q(\CPU_Xreg_value_a4[11][25] ),
    .CLK(clknet_8_183_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20350_ (.D(_00680_),
    .Q(\CPU_Xreg_value_a4[11][26] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20351_ (.D(_00681_),
    .Q(\CPU_Xreg_value_a4[11][27] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20352_ (.D(_00682_),
    .Q(\CPU_Xreg_value_a4[11][28] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20353_ (.D(_00683_),
    .Q(\CPU_Xreg_value_a4[11][29] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20354_ (.D(_00684_),
    .Q(\CPU_Xreg_value_a4[11][30] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20355_ (.D(_00685_),
    .Q(\CPU_Xreg_value_a4[11][31] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20356_ (.D(_00686_),
    .Q(\CPU_Xreg_value_a4[10][0] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20357_ (.D(_00687_),
    .Q(\CPU_Xreg_value_a4[10][1] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20358_ (.D(_00688_),
    .Q(\CPU_Xreg_value_a4[10][2] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20359_ (.D(_00689_),
    .Q(\CPU_Xreg_value_a4[10][3] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20360_ (.D(_00690_),
    .Q(\CPU_Xreg_value_a4[10][4] ),
    .CLK(clknet_8_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20361_ (.D(_00691_),
    .Q(\CPU_Xreg_value_a4[10][5] ),
    .CLK(clknet_8_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20362_ (.D(_00692_),
    .Q(\CPU_Xreg_value_a4[10][6] ),
    .CLK(clknet_8_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20363_ (.D(_00693_),
    .Q(\CPU_Xreg_value_a4[10][7] ),
    .CLK(clknet_8_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20364_ (.D(_00694_),
    .Q(\CPU_Xreg_value_a4[10][8] ),
    .CLK(clknet_8_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20365_ (.D(_00695_),
    .Q(\CPU_Xreg_value_a4[10][9] ),
    .CLK(clknet_8_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20366_ (.D(_00696_),
    .Q(\CPU_Xreg_value_a4[10][10] ),
    .CLK(clknet_8_19_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20367_ (.D(_00697_),
    .Q(\CPU_Xreg_value_a4[10][11] ),
    .CLK(clknet_8_26_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20368_ (.D(_00698_),
    .Q(\CPU_Xreg_value_a4[10][12] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20369_ (.D(_00699_),
    .Q(\CPU_Xreg_value_a4[10][13] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20370_ (.D(_00700_),
    .Q(\CPU_Xreg_value_a4[10][14] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20371_ (.D(_00701_),
    .Q(\CPU_Xreg_value_a4[10][15] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20372_ (.D(_00702_),
    .Q(\CPU_Xreg_value_a4[10][16] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20373_ (.D(_00703_),
    .Q(\CPU_Xreg_value_a4[10][17] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20374_ (.D(_00704_),
    .Q(\CPU_Xreg_value_a4[10][18] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20375_ (.D(_00705_),
    .Q(\CPU_Xreg_value_a4[10][19] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20376_ (.D(_00706_),
    .Q(\CPU_Xreg_value_a4[10][20] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20377_ (.D(_00707_),
    .Q(\CPU_Xreg_value_a4[10][21] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20378_ (.D(_00708_),
    .Q(\CPU_Xreg_value_a4[10][22] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20379_ (.D(_00709_),
    .Q(\CPU_Xreg_value_a4[10][23] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20380_ (.D(_00710_),
    .Q(\CPU_Xreg_value_a4[10][24] ),
    .CLK(clknet_8_183_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20381_ (.D(_00711_),
    .Q(\CPU_Xreg_value_a4[10][25] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20382_ (.D(_00712_),
    .Q(\CPU_Xreg_value_a4[10][26] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20383_ (.D(_00713_),
    .Q(\CPU_Xreg_value_a4[10][27] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20384_ (.D(_00714_),
    .Q(\CPU_Xreg_value_a4[10][28] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20385_ (.D(_00715_),
    .Q(\CPU_Xreg_value_a4[10][29] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20386_ (.D(_00716_),
    .Q(\CPU_Xreg_value_a4[10][30] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20387_ (.D(_00717_),
    .Q(\CPU_Xreg_value_a4[10][31] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20388_ (.D(_00718_),
    .Q(\CPU_Xreg_value_a4[9][0] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20389_ (.D(_00719_),
    .Q(\CPU_Xreg_value_a4[9][1] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20390_ (.D(_00720_),
    .Q(\CPU_Xreg_value_a4[9][2] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20391_ (.D(_00721_),
    .Q(\CPU_Xreg_value_a4[9][3] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20392_ (.D(_00722_),
    .Q(\CPU_Xreg_value_a4[9][4] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20393_ (.D(_00723_),
    .Q(\CPU_Xreg_value_a4[9][5] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20394_ (.D(_00724_),
    .Q(\CPU_Xreg_value_a4[9][6] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20395_ (.D(_00725_),
    .Q(\CPU_Xreg_value_a4[9][7] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20396_ (.D(_00726_),
    .Q(\CPU_Xreg_value_a4[9][8] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20397_ (.D(_00727_),
    .Q(\CPU_Xreg_value_a4[9][9] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20398_ (.D(_00728_),
    .Q(\CPU_Xreg_value_a4[9][10] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20399_ (.D(_00729_),
    .Q(\CPU_Xreg_value_a4[9][11] ),
    .CLK(clknet_8_16_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20400_ (.D(_00730_),
    .Q(\CPU_Xreg_value_a4[9][12] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20401_ (.D(_00731_),
    .Q(\CPU_Xreg_value_a4[9][13] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20402_ (.D(_00732_),
    .Q(\CPU_Xreg_value_a4[9][14] ),
    .CLK(clknet_8_29_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20403_ (.D(_00733_),
    .Q(\CPU_Xreg_value_a4[9][15] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20404_ (.D(_00734_),
    .Q(\CPU_Xreg_value_a4[9][16] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20405_ (.D(_00735_),
    .Q(\CPU_Xreg_value_a4[9][17] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20406_ (.D(_00736_),
    .Q(\CPU_Xreg_value_a4[9][18] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20407_ (.D(_00737_),
    .Q(\CPU_Xreg_value_a4[9][19] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20408_ (.D(_00738_),
    .Q(\CPU_Xreg_value_a4[9][20] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20409_ (.D(_00739_),
    .Q(\CPU_Xreg_value_a4[9][21] ),
    .CLK(clknet_8_158_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20410_ (.D(_00740_),
    .Q(\CPU_Xreg_value_a4[9][22] ),
    .CLK(clknet_8_180_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20411_ (.D(_00741_),
    .Q(\CPU_Xreg_value_a4[9][23] ),
    .CLK(clknet_8_177_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20412_ (.D(_00742_),
    .Q(\CPU_Xreg_value_a4[9][24] ),
    .CLK(clknet_8_182_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20413_ (.D(_00743_),
    .Q(\CPU_Xreg_value_a4[9][25] ),
    .CLK(clknet_8_188_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20414_ (.D(_00744_),
    .Q(\CPU_Xreg_value_a4[9][26] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20415_ (.D(_00745_),
    .Q(\CPU_Xreg_value_a4[9][27] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20416_ (.D(_00746_),
    .Q(\CPU_Xreg_value_a4[9][28] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20417_ (.D(_00747_),
    .Q(\CPU_Xreg_value_a4[9][29] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20418_ (.D(_00748_),
    .Q(\CPU_Xreg_value_a4[9][30] ),
    .CLK(clknet_8_147_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20419_ (.D(_00749_),
    .Q(\CPU_Xreg_value_a4[9][31] ),
    .CLK(clknet_8_150_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20420_ (.D(_00750_),
    .Q(\CPU_Xreg_value_a4[8][0] ),
    .CLK(clknet_8_145_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20421_ (.D(_00751_),
    .Q(\CPU_Xreg_value_a4[8][1] ),
    .CLK(clknet_8_144_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20422_ (.D(_00752_),
    .Q(\CPU_Xreg_value_a4[8][2] ),
    .CLK(clknet_8_58_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20423_ (.D(_00753_),
    .Q(\CPU_Xreg_value_a4[8][3] ),
    .CLK(clknet_8_147_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20424_ (.D(_00754_),
    .Q(\CPU_Xreg_value_a4[8][4] ),
    .CLK(clknet_8_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20425_ (.D(_00755_),
    .Q(\CPU_Xreg_value_a4[8][5] ),
    .CLK(clknet_8_39_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20426_ (.D(_00756_),
    .Q(\CPU_Xreg_value_a4[8][6] ),
    .CLK(clknet_8_37_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20427_ (.D(_00757_),
    .Q(\CPU_Xreg_value_a4[8][7] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20428_ (.D(_00758_),
    .Q(\CPU_Xreg_value_a4[8][8] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20429_ (.D(_00759_),
    .Q(\CPU_Xreg_value_a4[8][9] ),
    .CLK(clknet_8_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20430_ (.D(_00760_),
    .Q(\CPU_Xreg_value_a4[8][10] ),
    .CLK(clknet_8_18_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20431_ (.D(_00761_),
    .Q(\CPU_Xreg_value_a4[8][11] ),
    .CLK(clknet_8_7_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20432_ (.D(_00762_),
    .Q(\CPU_Xreg_value_a4[8][12] ),
    .CLK(clknet_8_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20433_ (.D(_00763_),
    .Q(\CPU_Xreg_value_a4[8][13] ),
    .CLK(clknet_8_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20434_ (.D(_00764_),
    .Q(\CPU_Xreg_value_a4[8][14] ),
    .CLK(clknet_8_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20435_ (.D(_00765_),
    .Q(\CPU_Xreg_value_a4[8][15] ),
    .CLK(clknet_8_49_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20436_ (.D(_00766_),
    .Q(\CPU_Xreg_value_a4[8][16] ),
    .CLK(clknet_8_48_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20437_ (.D(_00767_),
    .Q(\CPU_Xreg_value_a4[8][17] ),
    .CLK(clknet_8_50_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20438_ (.D(_00768_),
    .Q(\CPU_Xreg_value_a4[8][18] ),
    .CLK(clknet_8_56_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20439_ (.D(_00769_),
    .Q(\CPU_Xreg_value_a4[8][19] ),
    .CLK(clknet_8_155_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20440_ (.D(_00770_),
    .Q(\CPU_Xreg_value_a4[8][20] ),
    .CLK(clknet_8_155_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20441_ (.D(_00771_),
    .Q(\CPU_Xreg_value_a4[8][21] ),
    .CLK(clknet_8_155_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20442_ (.D(_00772_),
    .Q(\CPU_Xreg_value_a4[8][22] ),
    .CLK(clknet_8_177_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20443_ (.D(_00773_),
    .Q(\CPU_Xreg_value_a4[8][23] ),
    .CLK(clknet_8_177_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20444_ (.D(_00774_),
    .Q(\CPU_Xreg_value_a4[8][24] ),
    .CLK(clknet_8_179_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20445_ (.D(_00775_),
    .Q(\CPU_Xreg_value_a4[8][25] ),
    .CLK(clknet_8_190_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20446_ (.D(_00776_),
    .Q(\CPU_Xreg_value_a4[8][26] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20447_ (.D(_00777_),
    .Q(\CPU_Xreg_value_a4[8][27] ),
    .CLK(clknet_8_187_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20448_ (.D(_00778_),
    .Q(\CPU_Xreg_value_a4[8][28] ),
    .CLK(clknet_8_185_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20449_ (.D(_00779_),
    .Q(\CPU_Xreg_value_a4[8][29] ),
    .CLK(clknet_8_185_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20450_ (.D(_00780_),
    .Q(\CPU_Xreg_value_a4[8][30] ),
    .CLK(clknet_8_179_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20451_ (.D(_00781_),
    .Q(\CPU_Xreg_value_a4[8][31] ),
    .CLK(clknet_8_147_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20452_ (.D(_00782_),
    .Q(\CPU_Xreg_value_a4[7][0] ),
    .CLK(clknet_8_148_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20453_ (.D(_00783_),
    .Q(\CPU_Xreg_value_a4[7][1] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20454_ (.D(_00784_),
    .Q(\CPU_Xreg_value_a4[7][2] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20455_ (.D(_00785_),
    .Q(\CPU_Xreg_value_a4[7][3] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20456_ (.D(_00786_),
    .Q(\CPU_Xreg_value_a4[7][4] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20457_ (.D(_00787_),
    .Q(\CPU_Xreg_value_a4[7][5] ),
    .CLK(clknet_8_60_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20458_ (.D(_00788_),
    .Q(\CPU_Xreg_value_a4[7][6] ),
    .CLK(clknet_8_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20459_ (.D(_00789_),
    .Q(\CPU_Xreg_value_a4[7][7] ),
    .CLK(clknet_8_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20460_ (.D(_00790_),
    .Q(\CPU_Xreg_value_a4[7][8] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20461_ (.D(_00791_),
    .Q(\CPU_Xreg_value_a4[7][9] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20462_ (.D(_00792_),
    .Q(\CPU_Xreg_value_a4[7][10] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20463_ (.D(_00793_),
    .Q(\CPU_Xreg_value_a4[7][11] ),
    .CLK(clknet_8_17_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20464_ (.D(_00794_),
    .Q(\CPU_Xreg_value_a4[7][12] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20465_ (.D(_00795_),
    .Q(\CPU_Xreg_value_a4[7][13] ),
    .CLK(clknet_8_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20466_ (.D(_00796_),
    .Q(\CPU_Xreg_value_a4[7][14] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20467_ (.D(_00797_),
    .Q(\CPU_Xreg_value_a4[7][15] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20468_ (.D(_00798_),
    .Q(\CPU_Xreg_value_a4[7][16] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20469_ (.D(_00799_),
    .Q(\CPU_Xreg_value_a4[7][17] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20470_ (.D(_00800_),
    .Q(\CPU_Xreg_value_a4[7][18] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20471_ (.D(_00801_),
    .Q(\CPU_Xreg_value_a4[7][19] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20472_ (.D(_00802_),
    .Q(\CPU_Xreg_value_a4[7][20] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20473_ (.D(_00803_),
    .Q(\CPU_Xreg_value_a4[7][21] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20474_ (.D(_00804_),
    .Q(\CPU_Xreg_value_a4[7][22] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20475_ (.D(_00805_),
    .Q(\CPU_Xreg_value_a4[7][23] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20476_ (.D(_00806_),
    .Q(\CPU_Xreg_value_a4[7][24] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20477_ (.D(_00807_),
    .Q(\CPU_Xreg_value_a4[7][25] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20478_ (.D(_00808_),
    .Q(\CPU_Xreg_value_a4[7][26] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20479_ (.D(_00809_),
    .Q(\CPU_Xreg_value_a4[7][27] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20480_ (.D(_00810_),
    .Q(\CPU_Xreg_value_a4[7][28] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20481_ (.D(_00811_),
    .Q(\CPU_Xreg_value_a4[7][29] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20482_ (.D(_00812_),
    .Q(\CPU_Xreg_value_a4[7][30] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20483_ (.D(_00813_),
    .Q(\CPU_Xreg_value_a4[7][31] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20484_ (.D(_00814_),
    .Q(\CPU_Xreg_value_a4[6][0] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20485_ (.D(_00815_),
    .Q(\CPU_Xreg_value_a4[6][1] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20486_ (.D(_00816_),
    .Q(\CPU_Xreg_value_a4[6][2] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20487_ (.D(_00817_),
    .Q(\CPU_Xreg_value_a4[6][3] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20488_ (.D(_00818_),
    .Q(\CPU_Xreg_value_a4[6][4] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20489_ (.D(_00819_),
    .Q(\CPU_Xreg_value_a4[6][5] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20490_ (.D(_00820_),
    .Q(\CPU_Xreg_value_a4[6][6] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20491_ (.D(_00821_),
    .Q(\CPU_Xreg_value_a4[6][7] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20492_ (.D(_00822_),
    .Q(\CPU_Xreg_value_a4[6][8] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20493_ (.D(_00823_),
    .Q(\CPU_Xreg_value_a4[6][9] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20494_ (.D(_00824_),
    .Q(\CPU_Xreg_value_a4[6][10] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20495_ (.D(_00825_),
    .Q(\CPU_Xreg_value_a4[6][11] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20496_ (.D(_00826_),
    .Q(\CPU_Xreg_value_a4[6][12] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20497_ (.D(_00827_),
    .Q(\CPU_Xreg_value_a4[6][13] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20498_ (.D(_00828_),
    .Q(\CPU_Xreg_value_a4[6][14] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20499_ (.D(_00829_),
    .Q(\CPU_Xreg_value_a4[6][15] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20500_ (.D(_00830_),
    .Q(\CPU_Xreg_value_a4[6][16] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20501_ (.D(_00831_),
    .Q(\CPU_Xreg_value_a4[6][17] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20502_ (.D(_00832_),
    .Q(\CPU_Xreg_value_a4[6][18] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20503_ (.D(_00833_),
    .Q(\CPU_Xreg_value_a4[6][19] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20504_ (.D(_00834_),
    .Q(\CPU_Xreg_value_a4[6][20] ),
    .CLK(clknet_8_206_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20505_ (.D(_00835_),
    .Q(\CPU_Xreg_value_a4[6][21] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20506_ (.D(_00836_),
    .Q(\CPU_Xreg_value_a4[6][22] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20507_ (.D(_00837_),
    .Q(\CPU_Xreg_value_a4[6][23] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20508_ (.D(_00838_),
    .Q(\CPU_Xreg_value_a4[6][24] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20509_ (.D(_00839_),
    .Q(\CPU_Xreg_value_a4[6][25] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20510_ (.D(_00840_),
    .Q(\CPU_Xreg_value_a4[6][26] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20511_ (.D(_00841_),
    .Q(\CPU_Xreg_value_a4[6][27] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20512_ (.D(_00842_),
    .Q(\CPU_Xreg_value_a4[6][28] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20513_ (.D(_00843_),
    .Q(\CPU_Xreg_value_a4[6][29] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20514_ (.D(_00844_),
    .Q(\CPU_Xreg_value_a4[6][30] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20515_ (.D(_00845_),
    .Q(\CPU_Xreg_value_a4[6][31] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20516_ (.D(_00846_),
    .Q(\CPU_Xreg_value_a4[5][0] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20517_ (.D(_00847_),
    .Q(\CPU_Xreg_value_a4[5][1] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20518_ (.D(_00848_),
    .Q(\CPU_Xreg_value_a4[5][2] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20519_ (.D(_00849_),
    .Q(\CPU_Xreg_value_a4[5][3] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20520_ (.D(_00850_),
    .Q(\CPU_Xreg_value_a4[5][4] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20521_ (.D(_00851_),
    .Q(\CPU_Xreg_value_a4[5][5] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20522_ (.D(_00852_),
    .Q(\CPU_Xreg_value_a4[5][6] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20523_ (.D(_00853_),
    .Q(\CPU_Xreg_value_a4[5][7] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20524_ (.D(_00854_),
    .Q(\CPU_Xreg_value_a4[5][8] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20525_ (.D(_00855_),
    .Q(\CPU_Xreg_value_a4[5][9] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20526_ (.D(_00856_),
    .Q(\CPU_Xreg_value_a4[5][10] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20527_ (.D(_00857_),
    .Q(\CPU_Xreg_value_a4[5][11] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20528_ (.D(_00858_),
    .Q(\CPU_Xreg_value_a4[5][12] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20529_ (.D(_00859_),
    .Q(\CPU_Xreg_value_a4[5][13] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20530_ (.D(_00860_),
    .Q(\CPU_Xreg_value_a4[5][14] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20531_ (.D(_00861_),
    .Q(\CPU_Xreg_value_a4[5][15] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20532_ (.D(_00862_),
    .Q(\CPU_Xreg_value_a4[5][16] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20533_ (.D(_00863_),
    .Q(\CPU_Xreg_value_a4[5][17] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20534_ (.D(_00864_),
    .Q(\CPU_Xreg_value_a4[5][18] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20535_ (.D(_00865_),
    .Q(\CPU_Xreg_value_a4[5][19] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20536_ (.D(_00866_),
    .Q(\CPU_Xreg_value_a4[5][20] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20537_ (.D(_00867_),
    .Q(\CPU_Xreg_value_a4[5][21] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20538_ (.D(_00868_),
    .Q(\CPU_Xreg_value_a4[5][22] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20539_ (.D(_00869_),
    .Q(\CPU_Xreg_value_a4[5][23] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20540_ (.D(_00870_),
    .Q(\CPU_Xreg_value_a4[5][24] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20541_ (.D(_00871_),
    .Q(\CPU_Xreg_value_a4[5][25] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20542_ (.D(_00872_),
    .Q(\CPU_Xreg_value_a4[5][26] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20543_ (.D(_00873_),
    .Q(\CPU_Xreg_value_a4[5][27] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20544_ (.D(_00874_),
    .Q(\CPU_Xreg_value_a4[5][28] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20545_ (.D(_00875_),
    .Q(\CPU_Xreg_value_a4[5][29] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20546_ (.D(_00876_),
    .Q(\CPU_Xreg_value_a4[5][30] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20547_ (.D(_00877_),
    .Q(\CPU_Xreg_value_a4[5][31] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20548_ (.D(_00878_),
    .Q(\CPU_Xreg_value_a4[4][0] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20549_ (.D(_00879_),
    .Q(\CPU_Xreg_value_a4[4][1] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20550_ (.D(_00880_),
    .Q(\CPU_Xreg_value_a4[4][2] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20551_ (.D(_00881_),
    .Q(\CPU_Xreg_value_a4[4][3] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20552_ (.D(_00882_),
    .Q(\CPU_Xreg_value_a4[4][4] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20553_ (.D(_00883_),
    .Q(\CPU_Xreg_value_a4[4][5] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20554_ (.D(_00884_),
    .Q(\CPU_Xreg_value_a4[4][6] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20555_ (.D(_00885_),
    .Q(\CPU_Xreg_value_a4[4][7] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20556_ (.D(_00886_),
    .Q(\CPU_Xreg_value_a4[4][8] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20557_ (.D(_00887_),
    .Q(\CPU_Xreg_value_a4[4][9] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20558_ (.D(_00888_),
    .Q(\CPU_Xreg_value_a4[4][10] ),
    .CLK(clknet_8_23_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20559_ (.D(_00889_),
    .Q(\CPU_Xreg_value_a4[4][11] ),
    .CLK(clknet_8_28_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20560_ (.D(_00890_),
    .Q(\CPU_Xreg_value_a4[4][12] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20561_ (.D(_00891_),
    .Q(\CPU_Xreg_value_a4[4][13] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20562_ (.D(_00892_),
    .Q(\CPU_Xreg_value_a4[4][14] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20563_ (.D(_00893_),
    .Q(\CPU_Xreg_value_a4[4][15] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20564_ (.D(_00894_),
    .Q(\CPU_Xreg_value_a4[4][16] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20565_ (.D(_00895_),
    .Q(\CPU_Xreg_value_a4[4][17] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20566_ (.D(_00896_),
    .Q(\CPU_Xreg_value_a4[4][18] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20567_ (.D(_00897_),
    .Q(\CPU_Xreg_value_a4[4][19] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20568_ (.D(_00898_),
    .Q(\CPU_Xreg_value_a4[4][20] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20569_ (.D(_00899_),
    .Q(\CPU_Xreg_value_a4[4][21] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20570_ (.D(_00900_),
    .Q(\CPU_Xreg_value_a4[4][22] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20571_ (.D(_00901_),
    .Q(\CPU_Xreg_value_a4[4][23] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20572_ (.D(_00902_),
    .Q(\CPU_Xreg_value_a4[4][24] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20573_ (.D(_00903_),
    .Q(\CPU_Xreg_value_a4[4][25] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20574_ (.D(_00904_),
    .Q(\CPU_Xreg_value_a4[4][26] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20575_ (.D(_00905_),
    .Q(\CPU_Xreg_value_a4[4][27] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20576_ (.D(_00906_),
    .Q(\CPU_Xreg_value_a4[4][28] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20577_ (.D(_00907_),
    .Q(\CPU_Xreg_value_a4[4][29] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20578_ (.D(_00908_),
    .Q(\CPU_Xreg_value_a4[4][30] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20579_ (.D(_00909_),
    .Q(\CPU_Xreg_value_a4[4][31] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20580_ (.D(_00910_),
    .Q(\CPU_Xreg_value_a4[3][0] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20581_ (.D(_00911_),
    .Q(\CPU_Xreg_value_a4[3][1] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20582_ (.D(_00912_),
    .Q(\CPU_Xreg_value_a4[3][2] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20583_ (.D(_00913_),
    .Q(\CPU_Xreg_value_a4[3][3] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20584_ (.D(_00914_),
    .Q(\CPU_Xreg_value_a4[3][4] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20585_ (.D(_00915_),
    .Q(\CPU_Xreg_value_a4[3][5] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20586_ (.D(_00916_),
    .Q(\CPU_Xreg_value_a4[3][6] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20587_ (.D(_00917_),
    .Q(\CPU_Xreg_value_a4[3][7] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20588_ (.D(_00918_),
    .Q(\CPU_Xreg_value_a4[3][8] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20589_ (.D(_00919_),
    .Q(\CPU_Xreg_value_a4[3][9] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20590_ (.D(_00920_),
    .Q(\CPU_Xreg_value_a4[3][10] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20591_ (.D(_00921_),
    .Q(\CPU_Xreg_value_a4[3][11] ),
    .CLK(clknet_8_20_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20592_ (.D(_00922_),
    .Q(\CPU_Xreg_value_a4[3][12] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20593_ (.D(_00923_),
    .Q(\CPU_Xreg_value_a4[3][13] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20594_ (.D(_00924_),
    .Q(\CPU_Xreg_value_a4[3][14] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20595_ (.D(_00925_),
    .Q(\CPU_Xreg_value_a4[3][15] ),
    .CLK(clknet_8_22_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20596_ (.D(_00926_),
    .Q(\CPU_Xreg_value_a4[3][16] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20597_ (.D(_00927_),
    .Q(\CPU_Xreg_value_a4[3][17] ),
    .CLK(clknet_8_21_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20598_ (.D(_00928_),
    .Q(\CPU_Xreg_value_a4[3][18] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20599_ (.D(_00929_),
    .Q(\CPU_Xreg_value_a4[3][19] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20600_ (.D(_00930_),
    .Q(\CPU_Xreg_value_a4[3][20] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20601_ (.D(_00931_),
    .Q(\CPU_Xreg_value_a4[3][21] ),
    .CLK(clknet_8_202_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20602_ (.D(_00932_),
    .Q(\CPU_Xreg_value_a4[3][22] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20603_ (.D(_00933_),
    .Q(\CPU_Xreg_value_a4[3][23] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20604_ (.D(_00934_),
    .Q(\CPU_Xreg_value_a4[3][24] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20605_ (.D(_00935_),
    .Q(\CPU_Xreg_value_a4[3][25] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20606_ (.D(_00936_),
    .Q(\CPU_Xreg_value_a4[3][26] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20607_ (.D(_00937_),
    .Q(\CPU_Xreg_value_a4[3][27] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20608_ (.D(_00938_),
    .Q(\CPU_Xreg_value_a4[3][28] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20609_ (.D(_00939_),
    .Q(\CPU_Xreg_value_a4[3][29] ),
    .CLK(clknet_8_234_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20610_ (.D(_00940_),
    .Q(\CPU_Xreg_value_a4[3][30] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20611_ (.D(_00941_),
    .Q(\CPU_Xreg_value_a4[3][31] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20612_ (.D(_00942_),
    .Q(\CPU_Xreg_value_a4[2][0] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20613_ (.D(_00943_),
    .Q(\CPU_Xreg_value_a4[2][1] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20614_ (.D(_00944_),
    .Q(\CPU_Xreg_value_a4[2][2] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20615_ (.D(_00945_),
    .Q(\CPU_Xreg_value_a4[2][3] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20616_ (.D(_00946_),
    .Q(\CPU_Xreg_value_a4[2][4] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20617_ (.D(_00947_),
    .Q(\CPU_Xreg_value_a4[2][5] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20618_ (.D(_00948_),
    .Q(\CPU_Xreg_value_a4[2][6] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20619_ (.D(_00949_),
    .Q(\CPU_Xreg_value_a4[2][7] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20620_ (.D(_00950_),
    .Q(\CPU_Xreg_value_a4[2][8] ),
    .CLK(clknet_8_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20621_ (.D(_00951_),
    .Q(\CPU_Xreg_value_a4[2][9] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20622_ (.D(_00952_),
    .Q(\CPU_Xreg_value_a4[2][10] ),
    .CLK(clknet_8_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20623_ (.D(_00953_),
    .Q(\CPU_Xreg_value_a4[2][11] ),
    .CLK(clknet_8_25_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20624_ (.D(_00954_),
    .Q(\CPU_Xreg_value_a4[2][12] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20625_ (.D(_00955_),
    .Q(\CPU_Xreg_value_a4[2][13] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20626_ (.D(_00956_),
    .Q(\CPU_Xreg_value_a4[2][14] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20627_ (.D(_00957_),
    .Q(\CPU_Xreg_value_a4[2][15] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20628_ (.D(_00958_),
    .Q(\CPU_Xreg_value_a4[2][16] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20629_ (.D(_00959_),
    .Q(\CPU_Xreg_value_a4[2][17] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20630_ (.D(_00960_),
    .Q(\CPU_Xreg_value_a4[2][18] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20631_ (.D(_00961_),
    .Q(\CPU_Xreg_value_a4[2][19] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20632_ (.D(_00962_),
    .Q(\CPU_Xreg_value_a4[2][20] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20633_ (.D(_00963_),
    .Q(\CPU_Xreg_value_a4[2][21] ),
    .CLK(clknet_8_203_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20634_ (.D(_00964_),
    .Q(\CPU_Xreg_value_a4[2][22] ),
    .CLK(clknet_8_224_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20635_ (.D(_00965_),
    .Q(\CPU_Xreg_value_a4[2][23] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20636_ (.D(_00966_),
    .Q(\CPU_Xreg_value_a4[2][24] ),
    .CLK(clknet_8_226_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20637_ (.D(_00967_),
    .Q(\CPU_Xreg_value_a4[2][25] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20638_ (.D(_00968_),
    .Q(\CPU_Xreg_value_a4[2][26] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20639_ (.D(_00969_),
    .Q(\CPU_Xreg_value_a4[2][27] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20640_ (.D(_00970_),
    .Q(\CPU_Xreg_value_a4[2][28] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20641_ (.D(_00971_),
    .Q(\CPU_Xreg_value_a4[2][29] ),
    .CLK(clknet_8_232_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20642_ (.D(_00972_),
    .Q(\CPU_Xreg_value_a4[2][30] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20643_ (.D(_00973_),
    .Q(\CPU_Xreg_value_a4[2][31] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20644_ (.D(_00974_),
    .Q(\CPU_Xreg_value_a4[1][0] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20645_ (.D(_00975_),
    .Q(\CPU_Xreg_value_a4[1][1] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20646_ (.D(_00976_),
    .Q(\CPU_Xreg_value_a4[1][2] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20647_ (.D(_00977_),
    .Q(\CPU_Xreg_value_a4[1][3] ),
    .CLK(clknet_8_106_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20648_ (.D(_00978_),
    .Q(\CPU_Xreg_value_a4[1][4] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20649_ (.D(_00979_),
    .Q(\CPU_Xreg_value_a4[1][5] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20650_ (.D(_00980_),
    .Q(\CPU_Xreg_value_a4[1][6] ),
    .CLK(clknet_8_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20651_ (.D(_00981_),
    .Q(\CPU_Xreg_value_a4[1][7] ),
    .CLK(clknet_8_31_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20652_ (.D(_00982_),
    .Q(\CPU_Xreg_value_a4[1][8] ),
    .CLK(clknet_8_30_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20653_ (.D(_00983_),
    .Q(\CPU_Xreg_value_a4[1][9] ),
    .CLK(clknet_8_53_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20654_ (.D(_00984_),
    .Q(\CPU_Xreg_value_a4[1][10] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20655_ (.D(_00985_),
    .Q(\CPU_Xreg_value_a4[1][11] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20656_ (.D(_00986_),
    .Q(\CPU_Xreg_value_a4[1][12] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20657_ (.D(_00987_),
    .Q(\CPU_Xreg_value_a4[1][13] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20658_ (.D(_00988_),
    .Q(\CPU_Xreg_value_a4[1][14] ),
    .CLK(clknet_8_98_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20659_ (.D(_00989_),
    .Q(\CPU_Xreg_value_a4[1][15] ),
    .CLK(clknet_8_104_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20660_ (.D(_00990_),
    .Q(\CPU_Xreg_value_a4[1][16] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20661_ (.D(_00991_),
    .Q(\CPU_Xreg_value_a4[1][17] ),
    .CLK(clknet_8_195_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20662_ (.D(_00992_),
    .Q(\CPU_Xreg_value_a4[1][18] ),
    .CLK(clknet_8_201_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20663_ (.D(_00993_),
    .Q(\CPU_Xreg_value_a4[1][19] ),
    .CLK(clknet_8_204_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20664_ (.D(_00994_),
    .Q(\CPU_Xreg_value_a4[1][20] ),
    .CLK(clknet_8_206_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20665_ (.D(_00995_),
    .Q(\CPU_Xreg_value_a4[1][21] ),
    .CLK(clknet_8_206_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20666_ (.D(_00996_),
    .Q(\CPU_Xreg_value_a4[1][22] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20667_ (.D(_00997_),
    .Q(\CPU_Xreg_value_a4[1][23] ),
    .CLK(clknet_8_225_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20668_ (.D(_00998_),
    .Q(\CPU_Xreg_value_a4[1][24] ),
    .CLK(clknet_8_227_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20669_ (.D(_00999_),
    .Q(\CPU_Xreg_value_a4[1][25] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20670_ (.D(_01000_),
    .Q(\CPU_Xreg_value_a4[1][26] ),
    .CLK(clknet_8_235_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20671_ (.D(_01001_),
    .Q(\CPU_Xreg_value_a4[1][27] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20672_ (.D(_01002_),
    .Q(\CPU_Xreg_value_a4[1][28] ),
    .CLK(clknet_8_233_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20673_ (.D(_01003_),
    .Q(\CPU_Xreg_value_a4[1][29] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20674_ (.D(_01004_),
    .Q(\CPU_Xreg_value_a4[1][30] ),
    .CLK(clknet_8_194_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20675_ (.D(_01005_),
    .Q(\CPU_Xreg_value_a4[1][31] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20676_ (.D(_01006_),
    .Q(\CPU_Xreg_value_a4[0][0] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20677_ (.D(_01007_),
    .Q(\CPU_Xreg_value_a4[0][1] ),
    .CLK(clknet_8_149_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20678_ (.D(_01008_),
    .Q(\CPU_Xreg_value_a4[0][2] ),
    .CLK(clknet_8_192_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20679_ (.D(_01009_),
    .Q(\CPU_Xreg_value_a4[0][3] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20680_ (.D(_01010_),
    .Q(\CPU_Xreg_value_a4[0][4] ),
    .CLK(clknet_8_62_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20681_ (.D(_01011_),
    .Q(\CPU_Xreg_value_a4[0][5] ),
    .CLK(clknet_8_63_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20682_ (.D(_01012_),
    .Q(\CPU_Xreg_value_a4[0][6] ),
    .CLK(clknet_8_52_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20683_ (.D(_01013_),
    .Q(\CPU_Xreg_value_a4[0][7] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20684_ (.D(_01014_),
    .Q(\CPU_Xreg_value_a4[0][8] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20685_ (.D(_01015_),
    .Q(\CPU_Xreg_value_a4[0][9] ),
    .CLK(clknet_8_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20686_ (.D(_01016_),
    .Q(\CPU_Xreg_value_a4[0][10] ),
    .CLK(clknet_8_24_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20687_ (.D(_01017_),
    .Q(\CPU_Xreg_value_a4[0][11] ),
    .CLK(clknet_8_27_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20688_ (.D(_01018_),
    .Q(\CPU_Xreg_value_a4[0][12] ),
    .CLK(clknet_8_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20689_ (.D(_01019_),
    .Q(\CPU_Xreg_value_a4[0][13] ),
    .CLK(clknet_8_55_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20690_ (.D(_01020_),
    .Q(\CPU_Xreg_value_a4[0][14] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20691_ (.D(_01021_),
    .Q(\CPU_Xreg_value_a4[0][15] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20692_ (.D(_01022_),
    .Q(\CPU_Xreg_value_a4[0][16] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20693_ (.D(_01023_),
    .Q(\CPU_Xreg_value_a4[0][17] ),
    .CLK(clknet_8_61_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20694_ (.D(_01024_),
    .Q(\CPU_Xreg_value_a4[0][18] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20695_ (.D(_01025_),
    .Q(\CPU_Xreg_value_a4[0][19] ),
    .CLK(clknet_8_200_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20696_ (.D(_01026_),
    .Q(\CPU_Xreg_value_a4[0][20] ),
    .CLK(clknet_8_159_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20697_ (.D(_01027_),
    .Q(\CPU_Xreg_value_a4[0][21] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20698_ (.D(_01028_),
    .Q(\CPU_Xreg_value_a4[0][22] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20699_ (.D(_01029_),
    .Q(\CPU_Xreg_value_a4[0][23] ),
    .CLK(clknet_8_181_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20700_ (.D(_01030_),
    .Q(\CPU_Xreg_value_a4[0][24] ),
    .CLK(clknet_8_183_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20701_ (.D(_01031_),
    .Q(\CPU_Xreg_value_a4[0][25] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20702_ (.D(_01032_),
    .Q(\CPU_Xreg_value_a4[0][26] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20703_ (.D(_01033_),
    .Q(\CPU_Xreg_value_a4[0][27] ),
    .CLK(clknet_8_191_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20704_ (.D(_01034_),
    .Q(\CPU_Xreg_value_a4[0][28] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20705_ (.D(_01035_),
    .Q(\CPU_Xreg_value_a4[0][29] ),
    .CLK(clknet_8_189_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20706_ (.D(_01036_),
    .Q(\CPU_Xreg_value_a4[0][30] ),
    .CLK(clknet_8_157_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20707_ (.D(_01037_),
    .Q(\CPU_Xreg_value_a4[0][31] ),
    .CLK(clknet_8_151_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20708_ (.D(_01038_),
    .Q(\CPU_Dmem_value_a5[15][0] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20709_ (.D(_01039_),
    .Q(\CPU_Dmem_value_a5[15][1] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20710_ (.D(_01040_),
    .Q(\CPU_Dmem_value_a5[15][2] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20711_ (.D(_01041_),
    .Q(\CPU_Dmem_value_a5[15][3] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20712_ (.D(_01042_),
    .Q(\CPU_Dmem_value_a5[15][4] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20713_ (.D(_01043_),
    .Q(\CPU_Dmem_value_a5[15][5] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20714_ (.D(_01044_),
    .Q(\CPU_Dmem_value_a5[15][6] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20715_ (.D(_01045_),
    .Q(\CPU_Dmem_value_a5[15][7] ),
    .CLK(clknet_8_193_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20716_ (.D(_01046_),
    .Q(\CPU_Dmem_value_a5[15][8] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20717_ (.D(_01047_),
    .Q(\CPU_Dmem_value_a5[15][9] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20718_ (.D(_01048_),
    .Q(\CPU_Dmem_value_a5[15][10] ),
    .CLK(clknet_8_198_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20719_ (.D(_01049_),
    .Q(\CPU_Dmem_value_a5[15][11] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20720_ (.D(_01050_),
    .Q(\CPU_Dmem_value_a5[15][12] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20721_ (.D(_01051_),
    .Q(\CPU_Dmem_value_a5[15][13] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20722_ (.D(_01052_),
    .Q(\CPU_Dmem_value_a5[15][14] ),
    .CLK(clknet_8_199_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20723_ (.D(_01053_),
    .Q(\CPU_Dmem_value_a5[15][15] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20724_ (.D(_01054_),
    .Q(\CPU_Dmem_value_a5[15][16] ),
    .CLK(clknet_8_210_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20725_ (.D(_01055_),
    .Q(\CPU_Dmem_value_a5[15][17] ),
    .CLK(clknet_8_210_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20726_ (.D(_01056_),
    .Q(\CPU_Dmem_value_a5[15][18] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20727_ (.D(_01057_),
    .Q(\CPU_Dmem_value_a5[15][19] ),
    .CLK(clknet_8_220_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20728_ (.D(_01058_),
    .Q(\CPU_Dmem_value_a5[15][20] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20729_ (.D(_01059_),
    .Q(\CPU_Dmem_value_a5[15][21] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20730_ (.D(_01060_),
    .Q(\CPU_Dmem_value_a5[15][22] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20731_ (.D(_01061_),
    .Q(\CPU_Dmem_value_a5[15][23] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20732_ (.D(_01062_),
    .Q(\CPU_Dmem_value_a5[15][24] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20733_ (.D(_01063_),
    .Q(\CPU_Dmem_value_a5[15][25] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20734_ (.D(_01064_),
    .Q(\CPU_Dmem_value_a5[15][26] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20735_ (.D(_01065_),
    .Q(\CPU_Dmem_value_a5[15][27] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20736_ (.D(_01066_),
    .Q(\CPU_Dmem_value_a5[15][28] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20737_ (.D(_01067_),
    .Q(\CPU_Dmem_value_a5[15][29] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20738_ (.D(_01068_),
    .Q(\CPU_Dmem_value_a5[15][30] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20739_ (.D(_01069_),
    .Q(\CPU_Dmem_value_a5[15][31] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20740_ (.D(_01070_),
    .Q(\CPU_Dmem_value_a5[14][0] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20741_ (.D(_01071_),
    .Q(\CPU_Dmem_value_a5[14][1] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20742_ (.D(_01072_),
    .Q(\CPU_Dmem_value_a5[14][2] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20743_ (.D(_01073_),
    .Q(\CPU_Dmem_value_a5[14][3] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20744_ (.D(_01074_),
    .Q(\CPU_Dmem_value_a5[14][4] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20745_ (.D(_01075_),
    .Q(\CPU_Dmem_value_a5[14][5] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20746_ (.D(_01076_),
    .Q(\CPU_Dmem_value_a5[14][6] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20747_ (.D(_01077_),
    .Q(\CPU_Dmem_value_a5[14][7] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20748_ (.D(_01078_),
    .Q(\CPU_Dmem_value_a5[14][8] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20749_ (.D(_01079_),
    .Q(\CPU_Dmem_value_a5[14][9] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20750_ (.D(_01080_),
    .Q(\CPU_Dmem_value_a5[14][10] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20751_ (.D(_01081_),
    .Q(\CPU_Dmem_value_a5[14][11] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20752_ (.D(_01082_),
    .Q(\CPU_Dmem_value_a5[14][12] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20753_ (.D(_01083_),
    .Q(\CPU_Dmem_value_a5[14][13] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20754_ (.D(_01084_),
    .Q(\CPU_Dmem_value_a5[14][14] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20755_ (.D(_01085_),
    .Q(\CPU_Dmem_value_a5[14][15] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20756_ (.D(_01086_),
    .Q(\CPU_Dmem_value_a5[14][16] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20757_ (.D(_01087_),
    .Q(\CPU_Dmem_value_a5[14][17] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20758_ (.D(_01088_),
    .Q(\CPU_Dmem_value_a5[14][18] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20759_ (.D(_01089_),
    .Q(\CPU_Dmem_value_a5[14][19] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20760_ (.D(_01090_),
    .Q(\CPU_Dmem_value_a5[14][20] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20761_ (.D(_01091_),
    .Q(\CPU_Dmem_value_a5[14][21] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20762_ (.D(_01092_),
    .Q(\CPU_Dmem_value_a5[14][22] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20763_ (.D(_01093_),
    .Q(\CPU_Dmem_value_a5[14][23] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20764_ (.D(_01094_),
    .Q(\CPU_Dmem_value_a5[14][24] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20765_ (.D(_01095_),
    .Q(\CPU_Dmem_value_a5[14][25] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20766_ (.D(_01096_),
    .Q(\CPU_Dmem_value_a5[14][26] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20767_ (.D(_01097_),
    .Q(\CPU_Dmem_value_a5[14][27] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20768_ (.D(_01098_),
    .Q(\CPU_Dmem_value_a5[14][28] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20769_ (.D(_01099_),
    .Q(\CPU_Dmem_value_a5[14][29] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20770_ (.D(_01100_),
    .Q(\CPU_Dmem_value_a5[14][30] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20771_ (.D(_01101_),
    .Q(\CPU_Dmem_value_a5[14][31] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20772_ (.D(_01102_),
    .Q(\CPU_Dmem_value_a5[13][0] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20773_ (.D(_01103_),
    .Q(\CPU_Dmem_value_a5[13][1] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20774_ (.D(_01104_),
    .Q(\CPU_Dmem_value_a5[13][2] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20775_ (.D(_01105_),
    .Q(\CPU_Dmem_value_a5[13][3] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20776_ (.D(_01106_),
    .Q(\CPU_Dmem_value_a5[13][4] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20777_ (.D(_01107_),
    .Q(\CPU_Dmem_value_a5[13][5] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20778_ (.D(_01108_),
    .Q(\CPU_Dmem_value_a5[13][6] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20779_ (.D(_01109_),
    .Q(\CPU_Dmem_value_a5[13][7] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20780_ (.D(_01110_),
    .Q(\CPU_Dmem_value_a5[13][8] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20781_ (.D(_01111_),
    .Q(\CPU_Dmem_value_a5[13][9] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20782_ (.D(_01112_),
    .Q(\CPU_Dmem_value_a5[13][10] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20783_ (.D(_01113_),
    .Q(\CPU_Dmem_value_a5[13][11] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20784_ (.D(_01114_),
    .Q(\CPU_Dmem_value_a5[13][12] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20785_ (.D(_01115_),
    .Q(\CPU_Dmem_value_a5[13][13] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20786_ (.D(_01116_),
    .Q(\CPU_Dmem_value_a5[13][14] ),
    .CLK(clknet_8_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20787_ (.D(_01117_),
    .Q(\CPU_Dmem_value_a5[13][15] ),
    .CLK(clknet_8_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20788_ (.D(_01118_),
    .Q(\CPU_Dmem_value_a5[13][16] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20789_ (.D(_01119_),
    .Q(\CPU_Dmem_value_a5[13][17] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20790_ (.D(_01120_),
    .Q(\CPU_Dmem_value_a5[13][18] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20791_ (.D(_01121_),
    .Q(\CPU_Dmem_value_a5[13][19] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20792_ (.D(_01122_),
    .Q(\CPU_Dmem_value_a5[13][20] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20793_ (.D(_01123_),
    .Q(\CPU_Dmem_value_a5[13][21] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20794_ (.D(_01124_),
    .Q(\CPU_Dmem_value_a5[13][22] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20795_ (.D(_01125_),
    .Q(\CPU_Dmem_value_a5[13][23] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20796_ (.D(_01126_),
    .Q(\CPU_Dmem_value_a5[13][24] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20797_ (.D(_01127_),
    .Q(\CPU_Dmem_value_a5[13][25] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20798_ (.D(_01128_),
    .Q(\CPU_Dmem_value_a5[13][26] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20799_ (.D(_01129_),
    .Q(\CPU_Dmem_value_a5[13][27] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20800_ (.D(_01130_),
    .Q(\CPU_Dmem_value_a5[13][28] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20801_ (.D(_01131_),
    .Q(\CPU_Dmem_value_a5[13][29] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20802_ (.D(_01132_),
    .Q(\CPU_Dmem_value_a5[13][30] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20803_ (.D(_01133_),
    .Q(\CPU_Dmem_value_a5[13][31] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20804_ (.D(_01134_),
    .Q(\CPU_Dmem_value_a5[12][0] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20805_ (.D(_01135_),
    .Q(\CPU_Dmem_value_a5[12][1] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20806_ (.D(_01136_),
    .Q(\CPU_Dmem_value_a5[12][2] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20807_ (.D(_01137_),
    .Q(\CPU_Dmem_value_a5[12][3] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20808_ (.D(_01138_),
    .Q(\CPU_Dmem_value_a5[12][4] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20809_ (.D(_01139_),
    .Q(\CPU_Dmem_value_a5[12][5] ),
    .CLK(clknet_8_211_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20810_ (.D(_01140_),
    .Q(\CPU_Dmem_value_a5[12][6] ),
    .CLK(clknet_8_209_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20811_ (.D(_01141_),
    .Q(\CPU_Dmem_value_a5[12][7] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20812_ (.D(_01142_),
    .Q(\CPU_Dmem_value_a5[12][8] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20813_ (.D(_01143_),
    .Q(\CPU_Dmem_value_a5[12][9] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20814_ (.D(_01144_),
    .Q(\CPU_Dmem_value_a5[12][10] ),
    .CLK(clknet_8_196_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20815_ (.D(_01145_),
    .Q(\CPU_Dmem_value_a5[12][11] ),
    .CLK(clknet_8_197_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20816_ (.D(_01146_),
    .Q(\CPU_Dmem_value_a5[12][12] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20817_ (.D(_01147_),
    .Q(\CPU_Dmem_value_a5[12][13] ),
    .CLK(clknet_8_210_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20818_ (.D(_01148_),
    .Q(\CPU_Dmem_value_a5[12][14] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20819_ (.D(_01149_),
    .Q(\CPU_Dmem_value_a5[12][15] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20820_ (.D(_01150_),
    .Q(\CPU_Dmem_value_a5[12][16] ),
    .CLK(clknet_8_210_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20821_ (.D(_01151_),
    .Q(\CPU_Dmem_value_a5[12][17] ),
    .CLK(clknet_8_210_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20822_ (.D(_01152_),
    .Q(\CPU_Dmem_value_a5[12][18] ),
    .CLK(clknet_8_222_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20823_ (.D(_01153_),
    .Q(\CPU_Dmem_value_a5[12][19] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20824_ (.D(_01154_),
    .Q(\CPU_Dmem_value_a5[12][20] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20825_ (.D(_01155_),
    .Q(\CPU_Dmem_value_a5[12][21] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20826_ (.D(_01156_),
    .Q(\CPU_Dmem_value_a5[12][22] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20827_ (.D(_01157_),
    .Q(\CPU_Dmem_value_a5[12][23] ),
    .CLK(clknet_8_223_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20828_ (.D(_01158_),
    .Q(\CPU_Dmem_value_a5[12][24] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20829_ (.D(_01159_),
    .Q(\CPU_Dmem_value_a5[12][25] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20830_ (.D(_01160_),
    .Q(\CPU_Dmem_value_a5[12][26] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20831_ (.D(_01161_),
    .Q(\CPU_Dmem_value_a5[12][27] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20832_ (.D(_01162_),
    .Q(\CPU_Dmem_value_a5[12][28] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20833_ (.D(_01163_),
    .Q(\CPU_Dmem_value_a5[12][29] ),
    .CLK(clknet_8_221_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20834_ (.D(_01164_),
    .Q(\CPU_Dmem_value_a5[12][30] ),
    .CLK(clknet_8_215_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20835_ (.D(_01165_),
    .Q(\CPU_Dmem_value_a5[12][31] ),
    .CLK(clknet_8_214_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20836_ (.D(_01166_),
    .Q(\CPU_Dmem_value_a5[11][0] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20837_ (.D(_01167_),
    .Q(\CPU_Dmem_value_a5[11][1] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20838_ (.D(_01168_),
    .Q(\CPU_Dmem_value_a5[11][2] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20839_ (.D(_01169_),
    .Q(\CPU_Dmem_value_a5[11][3] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20840_ (.D(_01170_),
    .Q(\CPU_Dmem_value_a5[11][4] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20841_ (.D(_01171_),
    .Q(\CPU_Dmem_value_a5[11][5] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20842_ (.D(_01172_),
    .Q(\CPU_Dmem_value_a5[11][6] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20843_ (.D(_01173_),
    .Q(\CPU_Dmem_value_a5[11][7] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20844_ (.D(_01174_),
    .Q(\CPU_Dmem_value_a5[11][8] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20845_ (.D(_01175_),
    .Q(\CPU_Dmem_value_a5[11][9] ),
    .CLK(clknet_8_96_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20846_ (.D(_01176_),
    .Q(\CPU_Dmem_value_a5[11][10] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20847_ (.D(_01177_),
    .Q(\CPU_Dmem_value_a5[11][11] ),
    .CLK(clknet_8_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20848_ (.D(_01178_),
    .Q(\CPU_Dmem_value_a5[11][12] ),
    .CLK(clknet_8_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20849_ (.D(_01179_),
    .Q(\CPU_Dmem_value_a5[11][13] ),
    .CLK(clknet_8_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20850_ (.D(_01180_),
    .Q(\CPU_Dmem_value_a5[11][14] ),
    .CLK(clknet_8_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20851_ (.D(_01181_),
    .Q(\CPU_Dmem_value_a5[11][15] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20852_ (.D(_01182_),
    .Q(\CPU_Dmem_value_a5[11][16] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20853_ (.D(_01183_),
    .Q(\CPU_Dmem_value_a5[11][17] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20854_ (.D(_01184_),
    .Q(\CPU_Dmem_value_a5[11][18] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20855_ (.D(_01185_),
    .Q(\CPU_Dmem_value_a5[11][19] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20856_ (.D(_01186_),
    .Q(\CPU_Dmem_value_a5[11][20] ),
    .CLK(clknet_8_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20857_ (.D(_01187_),
    .Q(\CPU_Dmem_value_a5[11][21] ),
    .CLK(clknet_8_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20858_ (.D(_01188_),
    .Q(\CPU_Dmem_value_a5[11][22] ),
    .CLK(clknet_8_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20859_ (.D(_01189_),
    .Q(\CPU_Dmem_value_a5[11][23] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20860_ (.D(_01190_),
    .Q(\CPU_Dmem_value_a5[11][24] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20861_ (.D(_01191_),
    .Q(\CPU_Dmem_value_a5[11][25] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20862_ (.D(_01192_),
    .Q(\CPU_Dmem_value_a5[11][26] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20863_ (.D(_01193_),
    .Q(\CPU_Dmem_value_a5[11][27] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20864_ (.D(_01194_),
    .Q(\CPU_Dmem_value_a5[11][28] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20865_ (.D(_01195_),
    .Q(\CPU_Dmem_value_a5[11][29] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20866_ (.D(_01196_),
    .Q(\CPU_Dmem_value_a5[11][30] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20867_ (.D(_01197_),
    .Q(\CPU_Dmem_value_a5[11][31] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20868_ (.D(_01198_),
    .Q(\CPU_Dmem_value_a5[10][0] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20869_ (.D(_01199_),
    .Q(\CPU_Dmem_value_a5[10][1] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20870_ (.D(_01200_),
    .Q(\CPU_Dmem_value_a5[10][2] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20871_ (.D(_01201_),
    .Q(\CPU_Dmem_value_a5[10][3] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20872_ (.D(_01202_),
    .Q(\CPU_Dmem_value_a5[10][4] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20873_ (.D(_01203_),
    .Q(\CPU_Dmem_value_a5[10][5] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20874_ (.D(_01204_),
    .Q(\CPU_Dmem_value_a5[10][6] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20875_ (.D(_01205_),
    .Q(\CPU_Dmem_value_a5[10][7] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20876_ (.D(_01206_),
    .Q(\CPU_Dmem_value_a5[10][8] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20877_ (.D(_01207_),
    .Q(\CPU_Dmem_value_a5[10][9] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20878_ (.D(_01208_),
    .Q(\CPU_Dmem_value_a5[10][10] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20879_ (.D(_01209_),
    .Q(\CPU_Dmem_value_a5[10][11] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20880_ (.D(_01210_),
    .Q(\CPU_Dmem_value_a5[10][12] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20881_ (.D(_01211_),
    .Q(\CPU_Dmem_value_a5[10][13] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20882_ (.D(_01212_),
    .Q(\CPU_Dmem_value_a5[10][14] ),
    .CLK(clknet_8_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20883_ (.D(_01213_),
    .Q(\CPU_Dmem_value_a5[10][15] ),
    .CLK(clknet_8_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20884_ (.D(_01214_),
    .Q(\CPU_Dmem_value_a5[10][16] ),
    .CLK(clknet_8_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20885_ (.D(_01215_),
    .Q(\CPU_Dmem_value_a5[10][17] ),
    .CLK(clknet_8_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20886_ (.D(_01216_),
    .Q(\CPU_Dmem_value_a5[10][18] ),
    .CLK(clknet_8_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20887_ (.D(_01217_),
    .Q(\CPU_Dmem_value_a5[10][19] ),
    .CLK(clknet_8_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20888_ (.D(_01218_),
    .Q(\CPU_Dmem_value_a5[10][20] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20889_ (.D(_01219_),
    .Q(\CPU_Dmem_value_a5[10][21] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20890_ (.D(_01220_),
    .Q(\CPU_Dmem_value_a5[10][22] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20891_ (.D(_01221_),
    .Q(\CPU_Dmem_value_a5[10][23] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20892_ (.D(_01222_),
    .Q(\CPU_Dmem_value_a5[10][24] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20893_ (.D(_01223_),
    .Q(\CPU_Dmem_value_a5[10][25] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20894_ (.D(_01224_),
    .Q(\CPU_Dmem_value_a5[10][26] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20895_ (.D(_01225_),
    .Q(\CPU_Dmem_value_a5[10][27] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20896_ (.D(_01226_),
    .Q(\CPU_Dmem_value_a5[10][28] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20897_ (.D(_01227_),
    .Q(\CPU_Dmem_value_a5[10][29] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20898_ (.D(_01228_),
    .Q(\CPU_Dmem_value_a5[10][30] ),
    .CLK(clknet_8_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20899_ (.D(_01229_),
    .Q(\CPU_Dmem_value_a5[10][31] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20900_ (.D(_01230_),
    .Q(\CPU_Dmem_value_a5[9][0] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20901_ (.D(_01231_),
    .Q(\CPU_Dmem_value_a5[9][1] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20902_ (.D(_01232_),
    .Q(\CPU_Dmem_value_a5[9][2] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20903_ (.D(_01233_),
    .Q(\CPU_Dmem_value_a5[9][3] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20904_ (.D(_01234_),
    .Q(\CPU_Dmem_value_a5[9][4] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20905_ (.D(_01235_),
    .Q(\CPU_Dmem_value_a5[9][5] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20906_ (.D(_01236_),
    .Q(\CPU_Dmem_value_a5[9][6] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20907_ (.D(_01237_),
    .Q(\CPU_Dmem_value_a5[9][7] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20908_ (.D(_01238_),
    .Q(\CPU_Dmem_value_a5[9][8] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20909_ (.D(_01239_),
    .Q(\CPU_Dmem_value_a5[9][9] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20910_ (.D(_01240_),
    .Q(\CPU_Dmem_value_a5[9][10] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20911_ (.D(_01241_),
    .Q(\CPU_Dmem_value_a5[9][11] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20912_ (.D(_01242_),
    .Q(\CPU_Dmem_value_a5[9][12] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20913_ (.D(_01243_),
    .Q(\CPU_Dmem_value_a5[9][13] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20914_ (.D(_01244_),
    .Q(\CPU_Dmem_value_a5[9][14] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20915_ (.D(_01245_),
    .Q(\CPU_Dmem_value_a5[9][15] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20916_ (.D(_01246_),
    .Q(\CPU_Dmem_value_a5[9][16] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20917_ (.D(_01247_),
    .Q(\CPU_Dmem_value_a5[9][17] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20918_ (.D(_01248_),
    .Q(\CPU_Dmem_value_a5[9][18] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20919_ (.D(_01249_),
    .Q(\CPU_Dmem_value_a5[9][19] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20920_ (.D(_01250_),
    .Q(\CPU_Dmem_value_a5[9][20] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20921_ (.D(_01251_),
    .Q(\CPU_Dmem_value_a5[9][21] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20922_ (.D(_01252_),
    .Q(\CPU_Dmem_value_a5[9][22] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20923_ (.D(_01253_),
    .Q(\CPU_Dmem_value_a5[9][23] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20924_ (.D(_01254_),
    .Q(\CPU_Dmem_value_a5[9][24] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20925_ (.D(_01255_),
    .Q(\CPU_Dmem_value_a5[9][25] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20926_ (.D(_01256_),
    .Q(\CPU_Dmem_value_a5[9][26] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20927_ (.D(_01257_),
    .Q(\CPU_Dmem_value_a5[9][27] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20928_ (.D(_01258_),
    .Q(\CPU_Dmem_value_a5[9][28] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20929_ (.D(_01259_),
    .Q(\CPU_Dmem_value_a5[9][29] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20930_ (.D(_01260_),
    .Q(\CPU_Dmem_value_a5[9][30] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20931_ (.D(_01261_),
    .Q(\CPU_Dmem_value_a5[9][31] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20932_ (.D(_01262_),
    .Q(\CPU_Dmem_value_a5[8][0] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20933_ (.D(_01263_),
    .Q(\CPU_Dmem_value_a5[8][1] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20934_ (.D(_01264_),
    .Q(\CPU_Dmem_value_a5[8][2] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20935_ (.D(_01265_),
    .Q(\CPU_Dmem_value_a5[8][3] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20936_ (.D(_01266_),
    .Q(\CPU_Dmem_value_a5[8][4] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20937_ (.D(_01267_),
    .Q(\CPU_Dmem_value_a5[8][5] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20938_ (.D(_01268_),
    .Q(\CPU_Dmem_value_a5[8][6] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20939_ (.D(_01269_),
    .Q(\CPU_Dmem_value_a5[8][7] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20940_ (.D(_01270_),
    .Q(\CPU_Dmem_value_a5[8][8] ),
    .CLK(clknet_8_66_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20941_ (.D(_01271_),
    .Q(\CPU_Dmem_value_a5[8][9] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20942_ (.D(_01272_),
    .Q(\CPU_Dmem_value_a5[8][10] ),
    .CLK(clknet_8_67_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20943_ (.D(_01273_),
    .Q(\CPU_Dmem_value_a5[8][11] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20944_ (.D(_01274_),
    .Q(\CPU_Dmem_value_a5[8][12] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20945_ (.D(_01275_),
    .Q(\CPU_Dmem_value_a5[8][13] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20946_ (.D(_01276_),
    .Q(\CPU_Dmem_value_a5[8][14] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20947_ (.D(_01277_),
    .Q(\CPU_Dmem_value_a5[8][15] ),
    .CLK(clknet_8_70_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20948_ (.D(_01278_),
    .Q(\CPU_Dmem_value_a5[8][16] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20949_ (.D(_01279_),
    .Q(\CPU_Dmem_value_a5[8][17] ),
    .CLK(clknet_8_71_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20950_ (.D(_01280_),
    .Q(\CPU_Dmem_value_a5[8][18] ),
    .CLK(clknet_8_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20951_ (.D(_01281_),
    .Q(\CPU_Dmem_value_a5[8][19] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20952_ (.D(_01282_),
    .Q(\CPU_Dmem_value_a5[8][20] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20953_ (.D(_01283_),
    .Q(\CPU_Dmem_value_a5[8][21] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20954_ (.D(_01284_),
    .Q(\CPU_Dmem_value_a5[8][22] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20955_ (.D(_01285_),
    .Q(\CPU_Dmem_value_a5[8][23] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20956_ (.D(_01286_),
    .Q(\CPU_Dmem_value_a5[8][24] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20957_ (.D(_01287_),
    .Q(\CPU_Dmem_value_a5[8][25] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20958_ (.D(_01288_),
    .Q(\CPU_Dmem_value_a5[8][26] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20959_ (.D(_01289_),
    .Q(\CPU_Dmem_value_a5[8][27] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20960_ (.D(_01290_),
    .Q(\CPU_Dmem_value_a5[8][28] ),
    .CLK(clknet_8_87_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20961_ (.D(_01291_),
    .Q(\CPU_Dmem_value_a5[8][29] ),
    .CLK(clknet_8_86_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20962_ (.D(_01292_),
    .Q(\CPU_Dmem_value_a5[8][30] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20963_ (.D(_01293_),
    .Q(\CPU_Dmem_value_a5[8][31] ),
    .CLK(clknet_8_83_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20964_ (.D(_01294_),
    .Q(\CPU_Dmem_value_a5[7][0] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20965_ (.D(_01295_),
    .Q(\CPU_Dmem_value_a5[7][1] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20966_ (.D(_01296_),
    .Q(\CPU_Dmem_value_a5[7][2] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20967_ (.D(_01297_),
    .Q(\CPU_Dmem_value_a5[7][3] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20968_ (.D(_01298_),
    .Q(\CPU_Dmem_value_a5[7][4] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20969_ (.D(_01299_),
    .Q(\CPU_Dmem_value_a5[7][5] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20970_ (.D(_01300_),
    .Q(\CPU_Dmem_value_a5[7][6] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20971_ (.D(_01301_),
    .Q(\CPU_Dmem_value_a5[7][7] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20972_ (.D(_01302_),
    .Q(\CPU_Dmem_value_a5[7][8] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20973_ (.D(_01303_),
    .Q(\CPU_Dmem_value_a5[7][9] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20974_ (.D(_01304_),
    .Q(\CPU_Dmem_value_a5[7][10] ),
    .CLK(clknet_8_64_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20975_ (.D(_01305_),
    .Q(\CPU_Dmem_value_a5[7][11] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20976_ (.D(_01306_),
    .Q(\CPU_Dmem_value_a5[7][12] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20977_ (.D(_01307_),
    .Q(\CPU_Dmem_value_a5[7][13] ),
    .CLK(clknet_8_65_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20978_ (.D(_01308_),
    .Q(\CPU_Dmem_value_a5[7][14] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20979_ (.D(_01309_),
    .Q(\CPU_Dmem_value_a5[7][15] ),
    .CLK(clknet_8_68_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20980_ (.D(_01310_),
    .Q(\CPU_Dmem_value_a5[7][16] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20981_ (.D(_01311_),
    .Q(\CPU_Dmem_value_a5[7][17] ),
    .CLK(clknet_8_69_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20982_ (.D(_01312_),
    .Q(\CPU_Dmem_value_a5[7][18] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20983_ (.D(_01313_),
    .Q(\CPU_Dmem_value_a5[7][19] ),
    .CLK(clknet_8_80_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20984_ (.D(_01314_),
    .Q(\CPU_Dmem_value_a5[7][20] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20985_ (.D(_01315_),
    .Q(\CPU_Dmem_value_a5[7][21] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20986_ (.D(_01316_),
    .Q(\CPU_Dmem_value_a5[7][22] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20987_ (.D(_01317_),
    .Q(\CPU_Dmem_value_a5[7][23] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20988_ (.D(_01318_),
    .Q(\CPU_Dmem_value_a5[7][24] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20989_ (.D(_01319_),
    .Q(\CPU_Dmem_value_a5[7][25] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20990_ (.D(_01320_),
    .Q(\CPU_Dmem_value_a5[7][26] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20991_ (.D(_01321_),
    .Q(\CPU_Dmem_value_a5[7][27] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20992_ (.D(_01322_),
    .Q(\CPU_Dmem_value_a5[7][28] ),
    .CLK(clknet_8_85_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20993_ (.D(_01323_),
    .Q(\CPU_Dmem_value_a5[7][29] ),
    .CLK(clknet_8_84_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20994_ (.D(_01324_),
    .Q(\CPU_Dmem_value_a5[7][30] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20995_ (.D(_01325_),
    .Q(\CPU_Dmem_value_a5[7][31] ),
    .CLK(clknet_8_81_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20996_ (.D(_01326_),
    .Q(\CPU_Dmem_value_a5[6][0] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20997_ (.D(_01327_),
    .Q(\CPU_Dmem_value_a5[6][1] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20998_ (.D(_01328_),
    .Q(\CPU_Dmem_value_a5[6][2] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _20999_ (.D(_01329_),
    .Q(\CPU_Dmem_value_a5[6][3] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21000_ (.D(_01330_),
    .Q(\CPU_Dmem_value_a5[6][4] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21001_ (.D(_01331_),
    .Q(\CPU_Dmem_value_a5[6][5] ),
    .CLK(clknet_8_112_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21002_ (.D(_01332_),
    .Q(\CPU_Dmem_value_a5[6][6] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21003_ (.D(_01333_),
    .Q(\CPU_Dmem_value_a5[6][7] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21004_ (.D(_01334_),
    .Q(\CPU_Dmem_value_a5[6][8] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21005_ (.D(_01335_),
    .Q(\CPU_Dmem_value_a5[6][9] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21006_ (.D(_01336_),
    .Q(\CPU_Dmem_value_a5[6][10] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21007_ (.D(_01337_),
    .Q(\CPU_Dmem_value_a5[6][11] ),
    .CLK(clknet_8_97_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21008_ (.D(_01338_),
    .Q(\CPU_Dmem_value_a5[6][12] ),
    .CLK(clknet_8_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21009_ (.D(_01339_),
    .Q(\CPU_Dmem_value_a5[6][13] ),
    .CLK(clknet_8_100_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21010_ (.D(_01340_),
    .Q(\CPU_Dmem_value_a5[6][14] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21011_ (.D(_01341_),
    .Q(\CPU_Dmem_value_a5[6][15] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21012_ (.D(_01342_),
    .Q(\CPU_Dmem_value_a5[6][16] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21013_ (.D(_01343_),
    .Q(\CPU_Dmem_value_a5[6][17] ),
    .CLK(clknet_8_101_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21014_ (.D(_01344_),
    .Q(\CPU_Dmem_value_a5[6][18] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21015_ (.D(_01345_),
    .Q(\CPU_Dmem_value_a5[6][19] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21016_ (.D(_01346_),
    .Q(\CPU_Dmem_value_a5[6][20] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21017_ (.D(_01347_),
    .Q(\CPU_Dmem_value_a5[6][21] ),
    .CLK(clknet_8_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21018_ (.D(_01348_),
    .Q(\CPU_Dmem_value_a5[6][22] ),
    .CLK(clknet_8_118_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21019_ (.D(_01349_),
    .Q(\CPU_Dmem_value_a5[6][23] ),
    .CLK(clknet_8_116_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21020_ (.D(_01350_),
    .Q(\CPU_Dmem_value_a5[6][24] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21021_ (.D(_01351_),
    .Q(\CPU_Dmem_value_a5[6][25] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21022_ (.D(_01352_),
    .Q(\CPU_Dmem_value_a5[6][26] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21023_ (.D(_01353_),
    .Q(\CPU_Dmem_value_a5[6][27] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21024_ (.D(_01354_),
    .Q(\CPU_Dmem_value_a5[6][28] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21025_ (.D(_01355_),
    .Q(\CPU_Dmem_value_a5[6][29] ),
    .CLK(clknet_8_117_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21026_ (.D(_01356_),
    .Q(\CPU_Dmem_value_a5[6][30] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21027_ (.D(_01357_),
    .Q(\CPU_Dmem_value_a5[6][31] ),
    .CLK(clknet_8_113_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21028_ (.D(_01358_),
    .Q(\CPU_Dmem_value_a5[5][0] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21029_ (.D(_01359_),
    .Q(\CPU_Dmem_value_a5[5][1] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21030_ (.D(_01360_),
    .Q(\CPU_Dmem_value_a5[5][2] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21031_ (.D(_01361_),
    .Q(\CPU_Dmem_value_a5[5][3] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21032_ (.D(_01362_),
    .Q(\CPU_Dmem_value_a5[5][4] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21033_ (.D(_01363_),
    .Q(\CPU_Dmem_value_a5[5][5] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21034_ (.D(_01364_),
    .Q(\CPU_Dmem_value_a5[5][6] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21035_ (.D(_01365_),
    .Q(\CPU_Dmem_value_a5[5][7] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21036_ (.D(_01366_),
    .Q(\CPU_Dmem_value_a5[5][8] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21037_ (.D(_01367_),
    .Q(\CPU_Dmem_value_a5[5][9] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21038_ (.D(_01368_),
    .Q(\CPU_Dmem_value_a5[5][10] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21039_ (.D(_01369_),
    .Q(\CPU_Dmem_value_a5[5][11] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21040_ (.D(_01370_),
    .Q(\CPU_Dmem_value_a5[5][12] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21041_ (.D(_01371_),
    .Q(\CPU_Dmem_value_a5[5][13] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21042_ (.D(_01372_),
    .Q(\CPU_Dmem_value_a5[5][14] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21043_ (.D(_01373_),
    .Q(\CPU_Dmem_value_a5[5][15] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21044_ (.D(_01374_),
    .Q(\CPU_Dmem_value_a5[5][16] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21045_ (.D(_01375_),
    .Q(\CPU_Dmem_value_a5[5][17] ),
    .CLK(clknet_8_208_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21046_ (.D(_01376_),
    .Q(\CPU_Dmem_value_a5[5][18] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21047_ (.D(_01377_),
    .Q(\CPU_Dmem_value_a5[5][19] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21048_ (.D(_01378_),
    .Q(\CPU_Dmem_value_a5[5][20] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21049_ (.D(_01379_),
    .Q(\CPU_Dmem_value_a5[5][21] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21050_ (.D(_01380_),
    .Q(\CPU_Dmem_value_a5[5][22] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21051_ (.D(_01381_),
    .Q(\CPU_Dmem_value_a5[5][23] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21052_ (.D(_01382_),
    .Q(\CPU_Dmem_value_a5[5][24] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21053_ (.D(_01383_),
    .Q(\CPU_Dmem_value_a5[5][25] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21054_ (.D(_01384_),
    .Q(\CPU_Dmem_value_a5[5][26] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21055_ (.D(_01385_),
    .Q(\CPU_Dmem_value_a5[5][27] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21056_ (.D(_01386_),
    .Q(\CPU_Dmem_value_a5[5][28] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21057_ (.D(_01387_),
    .Q(\CPU_Dmem_value_a5[5][29] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21058_ (.D(_01388_),
    .Q(\CPU_Dmem_value_a5[5][30] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21059_ (.D(_01389_),
    .Q(\CPU_Dmem_value_a5[5][31] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21060_ (.D(_01390_),
    .Q(\CPU_Dmem_value_a5[4][0] ),
    .CLK(clknet_8_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21061_ (.D(_01391_),
    .Q(\CPU_Dmem_value_a5[4][1] ),
    .CLK(clknet_8_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21062_ (.D(_01392_),
    .Q(\CPU_Dmem_value_a5[4][2] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21063_ (.D(_01393_),
    .Q(\CPU_Dmem_value_a5[4][3] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21064_ (.D(_01394_),
    .Q(\CPU_Dmem_value_a5[4][4] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21065_ (.D(_01395_),
    .Q(\CPU_Dmem_value_a5[4][5] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21066_ (.D(_01396_),
    .Q(\CPU_Dmem_value_a5[4][6] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21067_ (.D(_01397_),
    .Q(\CPU_Dmem_value_a5[4][7] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21068_ (.D(_01398_),
    .Q(\CPU_Dmem_value_a5[4][8] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21069_ (.D(_01399_),
    .Q(\CPU_Dmem_value_a5[4][9] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21070_ (.D(_01400_),
    .Q(\CPU_Dmem_value_a5[4][10] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21071_ (.D(_01401_),
    .Q(\CPU_Dmem_value_a5[4][11] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21072_ (.D(_01402_),
    .Q(\CPU_Dmem_value_a5[4][12] ),
    .CLK(clknet_8_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21073_ (.D(_01403_),
    .Q(\CPU_Dmem_value_a5[4][13] ),
    .CLK(clknet_8_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21074_ (.D(_01404_),
    .Q(\CPU_Dmem_value_a5[4][14] ),
    .CLK(clknet_8_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21075_ (.D(_01405_),
    .Q(\CPU_Dmem_value_a5[4][15] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21076_ (.D(_01406_),
    .Q(\CPU_Dmem_value_a5[4][16] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21077_ (.D(_01407_),
    .Q(\CPU_Dmem_value_a5[4][17] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21078_ (.D(_01408_),
    .Q(\CPU_Dmem_value_a5[4][18] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21079_ (.D(_01409_),
    .Q(\CPU_Dmem_value_a5[4][19] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21080_ (.D(_01410_),
    .Q(\CPU_Dmem_value_a5[4][20] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21081_ (.D(_01411_),
    .Q(\CPU_Dmem_value_a5[4][21] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21082_ (.D(_01412_),
    .Q(\CPU_Dmem_value_a5[4][22] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21083_ (.D(_01413_),
    .Q(\CPU_Dmem_value_a5[4][23] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21084_ (.D(_01414_),
    .Q(\CPU_Dmem_value_a5[4][24] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21085_ (.D(_01415_),
    .Q(\CPU_Dmem_value_a5[4][25] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21086_ (.D(_01416_),
    .Q(\CPU_Dmem_value_a5[4][26] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21087_ (.D(_01417_),
    .Q(\CPU_Dmem_value_a5[4][27] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21088_ (.D(_01418_),
    .Q(\CPU_Dmem_value_a5[4][28] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21089_ (.D(_01419_),
    .Q(\CPU_Dmem_value_a5[4][29] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21090_ (.D(_01420_),
    .Q(\CPU_Dmem_value_a5[4][30] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21091_ (.D(_01421_),
    .Q(\CPU_Dmem_value_a5[4][31] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21092_ (.D(_01422_),
    .Q(\CPU_Dmem_value_a5[3][0] ),
    .CLK(clknet_8_82_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21093_ (.D(_01423_),
    .Q(\CPU_Dmem_value_a5[3][1] ),
    .CLK(clknet_8_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21094_ (.D(_01424_),
    .Q(\CPU_Dmem_value_a5[3][2] ),
    .CLK(clknet_8_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21095_ (.D(_01425_),
    .Q(\CPU_Dmem_value_a5[3][3] ),
    .CLK(clknet_8_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21096_ (.D(_01426_),
    .Q(\CPU_Dmem_value_a5[3][4] ),
    .CLK(clknet_8_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21097_ (.D(_01427_),
    .Q(\CPU_Dmem_value_a5[3][5] ),
    .CLK(clknet_8_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21098_ (.D(_01428_),
    .Q(\CPU_Dmem_value_a5[3][6] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21099_ (.D(_01429_),
    .Q(\CPU_Dmem_value_a5[3][7] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21100_ (.D(_01430_),
    .Q(\CPU_Dmem_value_a5[3][8] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21101_ (.D(_01431_),
    .Q(\CPU_Dmem_value_a5[3][9] ),
    .CLK(clknet_8_72_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21102_ (.D(_01432_),
    .Q(\CPU_Dmem_value_a5[3][10] ),
    .CLK(clknet_8_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21103_ (.D(_01433_),
    .Q(\CPU_Dmem_value_a5[3][11] ),
    .CLK(clknet_8_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21104_ (.D(_01434_),
    .Q(\CPU_Dmem_value_a5[3][12] ),
    .CLK(clknet_8_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21105_ (.D(_01435_),
    .Q(\CPU_Dmem_value_a5[3][13] ),
    .CLK(clknet_8_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21106_ (.D(_01436_),
    .Q(\CPU_Dmem_value_a5[3][14] ),
    .CLK(clknet_8_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21107_ (.D(_01437_),
    .Q(\CPU_Dmem_value_a5[3][15] ),
    .CLK(clknet_8_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21108_ (.D(_01438_),
    .Q(\CPU_Dmem_value_a5[3][16] ),
    .CLK(clknet_8_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21109_ (.D(_01439_),
    .Q(\CPU_Dmem_value_a5[3][17] ),
    .CLK(clknet_8_76_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21110_ (.D(_01440_),
    .Q(\CPU_Dmem_value_a5[3][18] ),
    .CLK(clknet_8_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21111_ (.D(_01441_),
    .Q(\CPU_Dmem_value_a5[3][19] ),
    .CLK(clknet_8_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21112_ (.D(_01442_),
    .Q(\CPU_Dmem_value_a5[3][20] ),
    .CLK(clknet_8_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21113_ (.D(_01443_),
    .Q(\CPU_Dmem_value_a5[3][21] ),
    .CLK(clknet_8_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21114_ (.D(_01444_),
    .Q(\CPU_Dmem_value_a5[3][22] ),
    .CLK(clknet_8_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21115_ (.D(_01445_),
    .Q(\CPU_Dmem_value_a5[3][23] ),
    .CLK(clknet_8_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21116_ (.D(_01446_),
    .Q(\CPU_Dmem_value_a5[3][24] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21117_ (.D(_01447_),
    .Q(\CPU_Dmem_value_a5[3][25] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21118_ (.D(_01448_),
    .Q(\CPU_Dmem_value_a5[3][26] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21119_ (.D(_01449_),
    .Q(\CPU_Dmem_value_a5[3][27] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21120_ (.D(_01450_),
    .Q(\CPU_Dmem_value_a5[3][28] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21121_ (.D(_01451_),
    .Q(\CPU_Dmem_value_a5[3][29] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21122_ (.D(_01452_),
    .Q(\CPU_Dmem_value_a5[3][30] ),
    .CLK(clknet_8_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21123_ (.D(_01453_),
    .Q(\CPU_Dmem_value_a5[3][31] ),
    .CLK(clknet_8_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21124_ (.D(_01454_),
    .Q(\CPU_Dmem_value_a5[2][0] ),
    .CLK(clknet_8_88_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21125_ (.D(_01455_),
    .Q(\CPU_Dmem_value_a5[2][1] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21126_ (.D(_01456_),
    .Q(\CPU_Dmem_value_a5[2][2] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21127_ (.D(_01457_),
    .Q(\CPU_Dmem_value_a5[2][3] ),
    .CLK(clknet_8_90_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21128_ (.D(_01458_),
    .Q(\CPU_Dmem_value_a5[2][4] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21129_ (.D(_01459_),
    .Q(\CPU_Dmem_value_a5[2][5] ),
    .CLK(clknet_8_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21130_ (.D(_01460_),
    .Q(\CPU_Dmem_value_a5[2][6] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21131_ (.D(_01461_),
    .Q(\CPU_Dmem_value_a5[2][7] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21132_ (.D(_01462_),
    .Q(\CPU_Dmem_value_a5[2][8] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21133_ (.D(_01463_),
    .Q(\CPU_Dmem_value_a5[2][9] ),
    .CLK(clknet_8_74_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21134_ (.D(_01464_),
    .Q(\CPU_Dmem_value_a5[2][10] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21135_ (.D(_01465_),
    .Q(\CPU_Dmem_value_a5[2][11] ),
    .CLK(clknet_8_73_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21136_ (.D(_01466_),
    .Q(\CPU_Dmem_value_a5[2][12] ),
    .CLK(clknet_8_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21137_ (.D(_01467_),
    .Q(\CPU_Dmem_value_a5[2][13] ),
    .CLK(clknet_8_75_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21138_ (.D(_01468_),
    .Q(\CPU_Dmem_value_a5[2][14] ),
    .CLK(clknet_8_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21139_ (.D(_01469_),
    .Q(\CPU_Dmem_value_a5[2][15] ),
    .CLK(clknet_8_78_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21140_ (.D(_01470_),
    .Q(\CPU_Dmem_value_a5[2][16] ),
    .CLK(clknet_8_77_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21141_ (.D(_01471_),
    .Q(\CPU_Dmem_value_a5[2][17] ),
    .CLK(clknet_8_79_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21142_ (.D(_01472_),
    .Q(\CPU_Dmem_value_a5[2][18] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21143_ (.D(_01473_),
    .Q(\CPU_Dmem_value_a5[2][19] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21144_ (.D(_01474_),
    .Q(\CPU_Dmem_value_a5[2][20] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21145_ (.D(_01475_),
    .Q(\CPU_Dmem_value_a5[2][21] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21146_ (.D(_01476_),
    .Q(\CPU_Dmem_value_a5[2][22] ),
    .CLK(clknet_8_92_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21147_ (.D(_01477_),
    .Q(\CPU_Dmem_value_a5[2][23] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21148_ (.D(_01478_),
    .Q(\CPU_Dmem_value_a5[2][24] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21149_ (.D(_01479_),
    .Q(\CPU_Dmem_value_a5[2][25] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21150_ (.D(_01480_),
    .Q(\CPU_Dmem_value_a5[2][26] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21151_ (.D(_01481_),
    .Q(\CPU_Dmem_value_a5[2][27] ),
    .CLK(clknet_8_95_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21152_ (.D(_01482_),
    .Q(\CPU_Dmem_value_a5[2][28] ),
    .CLK(clknet_8_94_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21153_ (.D(_01483_),
    .Q(\CPU_Dmem_value_a5[2][29] ),
    .CLK(clknet_8_93_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21154_ (.D(_01484_),
    .Q(\CPU_Dmem_value_a5[2][30] ),
    .CLK(clknet_8_91_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21155_ (.D(_01485_),
    .Q(\CPU_Dmem_value_a5[2][31] ),
    .CLK(clknet_8_89_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21156_ (.D(_01486_),
    .Q(\CPU_Dmem_value_a5[1][0] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21157_ (.D(_01487_),
    .Q(\CPU_Dmem_value_a5[1][1] ),
    .CLK(clknet_8_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21158_ (.D(_01488_),
    .Q(\CPU_Dmem_value_a5[1][2] ),
    .CLK(clknet_8_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21159_ (.D(_01489_),
    .Q(\CPU_Dmem_value_a5[1][3] ),
    .CLK(clknet_8_115_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21160_ (.D(_01490_),
    .Q(\CPU_Dmem_value_a5[1][4] ),
    .CLK(clknet_8_114_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21161_ (.D(_01491_),
    .Q(\CPU_Dmem_value_a5[1][5] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21162_ (.D(_01492_),
    .Q(\CPU_Dmem_value_a5[1][6] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21163_ (.D(_01493_),
    .Q(\CPU_Dmem_value_a5[1][7] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21164_ (.D(_01494_),
    .Q(\CPU_Dmem_value_a5[1][8] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21165_ (.D(_01495_),
    .Q(\CPU_Dmem_value_a5[1][9] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21166_ (.D(_01496_),
    .Q(\CPU_Dmem_value_a5[1][10] ),
    .CLK(clknet_8_99_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21167_ (.D(_01497_),
    .Q(\CPU_Dmem_value_a5[1][11] ),
    .CLK(clknet_8_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21168_ (.D(_01498_),
    .Q(\CPU_Dmem_value_a5[1][12] ),
    .CLK(clknet_8_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21169_ (.D(_01499_),
    .Q(\CPU_Dmem_value_a5[1][13] ),
    .CLK(clknet_8_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21170_ (.D(_01500_),
    .Q(\CPU_Dmem_value_a5[1][14] ),
    .CLK(clknet_8_102_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21171_ (.D(_01501_),
    .Q(\CPU_Dmem_value_a5[1][15] ),
    .CLK(clknet_8_103_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21172_ (.D(_01502_),
    .Q(\CPU_Dmem_value_a5[1][16] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21173_ (.D(_01503_),
    .Q(\CPU_Dmem_value_a5[1][17] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21174_ (.D(_01504_),
    .Q(\CPU_Dmem_value_a5[1][18] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21175_ (.D(_01505_),
    .Q(\CPU_Dmem_value_a5[1][19] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21176_ (.D(_01506_),
    .Q(\CPU_Dmem_value_a5[1][20] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21177_ (.D(_01507_),
    .Q(\CPU_Dmem_value_a5[1][21] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21178_ (.D(_01508_),
    .Q(\CPU_Dmem_value_a5[1][22] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21179_ (.D(_01509_),
    .Q(\CPU_Dmem_value_a5[1][23] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21180_ (.D(_01510_),
    .Q(\CPU_Dmem_value_a5[1][24] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21181_ (.D(_01511_),
    .Q(\CPU_Dmem_value_a5[1][25] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21182_ (.D(_01512_),
    .Q(\CPU_Dmem_value_a5[1][26] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21183_ (.D(_01513_),
    .Q(\CPU_Dmem_value_a5[1][27] ),
    .CLK(clknet_8_119_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21184_ (.D(_01514_),
    .Q(\CPU_Dmem_value_a5[1][28] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21185_ (.D(_01515_),
    .Q(\CPU_Dmem_value_a5[1][29] ),
    .CLK(clknet_8_125_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21186_ (.D(_01516_),
    .Q(\CPU_Dmem_value_a5[1][30] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21187_ (.D(_01517_),
    .Q(\CPU_Dmem_value_a5[1][31] ),
    .CLK(clknet_8_124_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21188_ (.D(_01518_),
    .Q(\CPU_Dmem_value_a5[0][0] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21189_ (.D(_01519_),
    .Q(\CPU_Dmem_value_a5[0][1] ),
    .CLK(clknet_8_121_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21190_ (.D(_01520_),
    .Q(\CPU_Dmem_value_a5[0][2] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21191_ (.D(_01521_),
    .Q(\CPU_Dmem_value_a5[0][3] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21192_ (.D(_01522_),
    .Q(\CPU_Dmem_value_a5[0][4] ),
    .CLK(clknet_8_120_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21193_ (.D(_01523_),
    .Q(\CPU_Dmem_value_a5[0][5] ),
    .CLK(clknet_8_109_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21194_ (.D(_01524_),
    .Q(\CPU_Dmem_value_a5[0][6] ),
    .CLK(clknet_8_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21195_ (.D(_01525_),
    .Q(\CPU_Dmem_value_a5[0][7] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21196_ (.D(_01526_),
    .Q(\CPU_Dmem_value_a5[0][8] ),
    .CLK(clknet_8_105_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21197_ (.D(_01527_),
    .Q(\CPU_Dmem_value_a5[0][9] ),
    .CLK(clknet_8_107_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21198_ (.D(_01528_),
    .Q(\CPU_Dmem_value_a5[0][10] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21199_ (.D(_01529_),
    .Q(\CPU_Dmem_value_a5[0][11] ),
    .CLK(clknet_8_110_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21200_ (.D(_01530_),
    .Q(\CPU_Dmem_value_a5[0][12] ),
    .CLK(clknet_8_108_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21201_ (.D(_01531_),
    .Q(\CPU_Dmem_value_a5[0][13] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21202_ (.D(_01532_),
    .Q(\CPU_Dmem_value_a5[0][14] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21203_ (.D(_01533_),
    .Q(\CPU_Dmem_value_a5[0][15] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21204_ (.D(_01534_),
    .Q(\CPU_Dmem_value_a5[0][16] ),
    .CLK(clknet_8_111_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21205_ (.D(_01535_),
    .Q(\CPU_Dmem_value_a5[0][17] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21206_ (.D(_01536_),
    .Q(\CPU_Dmem_value_a5[0][18] ),
    .CLK(clknet_8_122_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21207_ (.D(_01537_),
    .Q(\CPU_Dmem_value_a5[0][19] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21208_ (.D(_01538_),
    .Q(\CPU_Dmem_value_a5[0][20] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21209_ (.D(_01539_),
    .Q(\CPU_Dmem_value_a5[0][21] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21210_ (.D(_01540_),
    .Q(\CPU_Dmem_value_a5[0][22] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21211_ (.D(_01541_),
    .Q(\CPU_Dmem_value_a5[0][23] ),
    .CLK(clknet_8_213_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21212_ (.D(_01542_),
    .Q(\CPU_Dmem_value_a5[0][24] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21213_ (.D(_01543_),
    .Q(\CPU_Dmem_value_a5[0][25] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21214_ (.D(_01544_),
    .Q(\CPU_Dmem_value_a5[0][26] ),
    .CLK(clknet_8_212_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21215_ (.D(_01545_),
    .Q(\CPU_Dmem_value_a5[0][27] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21216_ (.D(_01546_),
    .Q(\CPU_Dmem_value_a5[0][28] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21217_ (.D(_01547_),
    .Q(\CPU_Dmem_value_a5[0][29] ),
    .CLK(clknet_8_127_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21218_ (.D(_01548_),
    .Q(\CPU_Dmem_value_a5[0][30] ),
    .CLK(clknet_8_126_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _21219_ (.D(_01549_),
    .Q(\CPU_Dmem_value_a5[0][31] ),
    .CLK(clknet_8_123_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_2_0_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_1_clk (.A(clknet_2_1_0_clk),
    .X(clknet_2_1_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_1_clk (.A(clknet_2_2_0_clk),
    .X(clknet_2_2_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_1_clk (.A(clknet_2_3_0_clk),
    .X(clknet_2_3_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_0_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_1_0_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_2_0_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_3_0_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_4_0_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_5_0_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_6_0_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_7_0_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_8_0_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_9_0_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_10_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_11_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_12_0_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_13_0_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_14_0_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_15_0_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_16_0_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_17_0_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_18_0_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_19_0_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_20_0_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_21_0_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_22_0_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_23_0_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_24_0_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_25_0_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_26_0_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_27_0_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_28_0_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_29_0_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_30_0_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_31_0_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_32_0_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_33_0_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_34_0_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_35_0_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_36_0_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_37_0_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_38_0_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_39_0_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_40_0_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_41_0_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_42_0_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_43_0_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_44_0_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_45_0_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_46_0_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_47_0_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_48_0_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_49_0_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_50_0_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_51_0_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_52_0_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_53_0_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_54_0_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_55_0_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_56_0_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_57_0_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_58_0_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_59_0_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_60_0_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_61_0_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_62_0_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_6_63_0_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_0_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_7_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_1_0_clk (.A(clknet_6_0_0_clk),
    .X(clknet_7_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_2_0_clk (.A(clknet_6_1_0_clk),
    .X(clknet_7_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_3_0_clk (.A(clknet_6_1_0_clk),
    .X(clknet_7_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_4_0_clk (.A(clknet_6_2_0_clk),
    .X(clknet_7_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_5_0_clk (.A(clknet_6_2_0_clk),
    .X(clknet_7_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_6_0_clk (.A(clknet_6_3_0_clk),
    .X(clknet_7_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_7_0_clk (.A(clknet_6_3_0_clk),
    .X(clknet_7_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_8_0_clk (.A(clknet_6_4_0_clk),
    .X(clknet_7_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_9_0_clk (.A(clknet_6_4_0_clk),
    .X(clknet_7_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_10_0_clk (.A(clknet_6_5_0_clk),
    .X(clknet_7_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_11_0_clk (.A(clknet_6_5_0_clk),
    .X(clknet_7_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_12_0_clk (.A(clknet_6_6_0_clk),
    .X(clknet_7_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_13_0_clk (.A(clknet_6_6_0_clk),
    .X(clknet_7_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_14_0_clk (.A(clknet_6_7_0_clk),
    .X(clknet_7_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_15_0_clk (.A(clknet_6_7_0_clk),
    .X(clknet_7_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_16_0_clk (.A(clknet_6_8_0_clk),
    .X(clknet_7_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_17_0_clk (.A(clknet_6_8_0_clk),
    .X(clknet_7_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_18_0_clk (.A(clknet_6_9_0_clk),
    .X(clknet_7_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_19_0_clk (.A(clknet_6_9_0_clk),
    .X(clknet_7_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_20_0_clk (.A(clknet_6_10_0_clk),
    .X(clknet_7_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_21_0_clk (.A(clknet_6_10_0_clk),
    .X(clknet_7_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_22_0_clk (.A(clknet_6_11_0_clk),
    .X(clknet_7_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_23_0_clk (.A(clknet_6_11_0_clk),
    .X(clknet_7_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_24_0_clk (.A(clknet_6_12_0_clk),
    .X(clknet_7_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_25_0_clk (.A(clknet_6_12_0_clk),
    .X(clknet_7_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_26_0_clk (.A(clknet_6_13_0_clk),
    .X(clknet_7_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_27_0_clk (.A(clknet_6_13_0_clk),
    .X(clknet_7_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_28_0_clk (.A(clknet_6_14_0_clk),
    .X(clknet_7_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_29_0_clk (.A(clknet_6_14_0_clk),
    .X(clknet_7_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_30_0_clk (.A(clknet_6_15_0_clk),
    .X(clknet_7_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_31_0_clk (.A(clknet_6_15_0_clk),
    .X(clknet_7_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_32_0_clk (.A(clknet_6_16_0_clk),
    .X(clknet_7_32_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_33_0_clk (.A(clknet_6_16_0_clk),
    .X(clknet_7_33_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_34_0_clk (.A(clknet_6_17_0_clk),
    .X(clknet_7_34_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_35_0_clk (.A(clknet_6_17_0_clk),
    .X(clknet_7_35_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_36_0_clk (.A(clknet_6_18_0_clk),
    .X(clknet_7_36_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_37_0_clk (.A(clknet_6_18_0_clk),
    .X(clknet_7_37_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_38_0_clk (.A(clknet_6_19_0_clk),
    .X(clknet_7_38_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_39_0_clk (.A(clknet_6_19_0_clk),
    .X(clknet_7_39_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_40_0_clk (.A(clknet_6_20_0_clk),
    .X(clknet_7_40_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_41_0_clk (.A(clknet_6_20_0_clk),
    .X(clknet_7_41_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_42_0_clk (.A(clknet_6_21_0_clk),
    .X(clknet_7_42_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_43_0_clk (.A(clknet_6_21_0_clk),
    .X(clknet_7_43_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_44_0_clk (.A(clknet_6_22_0_clk),
    .X(clknet_7_44_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_45_0_clk (.A(clknet_6_22_0_clk),
    .X(clknet_7_45_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_46_0_clk (.A(clknet_6_23_0_clk),
    .X(clknet_7_46_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_47_0_clk (.A(clknet_6_23_0_clk),
    .X(clknet_7_47_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_48_0_clk (.A(clknet_6_24_0_clk),
    .X(clknet_7_48_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_49_0_clk (.A(clknet_6_24_0_clk),
    .X(clknet_7_49_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_50_0_clk (.A(clknet_6_25_0_clk),
    .X(clknet_7_50_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_51_0_clk (.A(clknet_6_25_0_clk),
    .X(clknet_7_51_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_52_0_clk (.A(clknet_6_26_0_clk),
    .X(clknet_7_52_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_53_0_clk (.A(clknet_6_26_0_clk),
    .X(clknet_7_53_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_54_0_clk (.A(clknet_6_27_0_clk),
    .X(clknet_7_54_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_55_0_clk (.A(clknet_6_27_0_clk),
    .X(clknet_7_55_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_56_0_clk (.A(clknet_6_28_0_clk),
    .X(clknet_7_56_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_57_0_clk (.A(clknet_6_28_0_clk),
    .X(clknet_7_57_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_58_0_clk (.A(clknet_6_29_0_clk),
    .X(clknet_7_58_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_59_0_clk (.A(clknet_6_29_0_clk),
    .X(clknet_7_59_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_60_0_clk (.A(clknet_6_30_0_clk),
    .X(clknet_7_60_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_61_0_clk (.A(clknet_6_30_0_clk),
    .X(clknet_7_61_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_62_0_clk (.A(clknet_6_31_0_clk),
    .X(clknet_7_62_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_63_0_clk (.A(clknet_6_31_0_clk),
    .X(clknet_7_63_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_64_0_clk (.A(clknet_6_32_0_clk),
    .X(clknet_7_64_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_65_0_clk (.A(clknet_6_32_0_clk),
    .X(clknet_7_65_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_66_0_clk (.A(clknet_6_33_0_clk),
    .X(clknet_7_66_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_67_0_clk (.A(clknet_6_33_0_clk),
    .X(clknet_7_67_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_68_0_clk (.A(clknet_6_34_0_clk),
    .X(clknet_7_68_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_69_0_clk (.A(clknet_6_34_0_clk),
    .X(clknet_7_69_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_70_0_clk (.A(clknet_6_35_0_clk),
    .X(clknet_7_70_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_71_0_clk (.A(clknet_6_35_0_clk),
    .X(clknet_7_71_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_72_0_clk (.A(clknet_6_36_0_clk),
    .X(clknet_7_72_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_73_0_clk (.A(clknet_6_36_0_clk),
    .X(clknet_7_73_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_74_0_clk (.A(clknet_6_37_0_clk),
    .X(clknet_7_74_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_75_0_clk (.A(clknet_6_37_0_clk),
    .X(clknet_7_75_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_76_0_clk (.A(clknet_6_38_0_clk),
    .X(clknet_7_76_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_77_0_clk (.A(clknet_6_38_0_clk),
    .X(clknet_7_77_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_78_0_clk (.A(clknet_6_39_0_clk),
    .X(clknet_7_78_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_79_0_clk (.A(clknet_6_39_0_clk),
    .X(clknet_7_79_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_80_0_clk (.A(clknet_6_40_0_clk),
    .X(clknet_7_80_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_81_0_clk (.A(clknet_6_40_0_clk),
    .X(clknet_7_81_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_82_0_clk (.A(clknet_6_41_0_clk),
    .X(clknet_7_82_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_83_0_clk (.A(clknet_6_41_0_clk),
    .X(clknet_7_83_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_84_0_clk (.A(clknet_6_42_0_clk),
    .X(clknet_7_84_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_85_0_clk (.A(clknet_6_42_0_clk),
    .X(clknet_7_85_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_86_0_clk (.A(clknet_6_43_0_clk),
    .X(clknet_7_86_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_87_0_clk (.A(clknet_6_43_0_clk),
    .X(clknet_7_87_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_88_0_clk (.A(clknet_6_44_0_clk),
    .X(clknet_7_88_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_89_0_clk (.A(clknet_6_44_0_clk),
    .X(clknet_7_89_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_90_0_clk (.A(clknet_6_45_0_clk),
    .X(clknet_7_90_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_91_0_clk (.A(clknet_6_45_0_clk),
    .X(clknet_7_91_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_92_0_clk (.A(clknet_6_46_0_clk),
    .X(clknet_7_92_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_93_0_clk (.A(clknet_6_46_0_clk),
    .X(clknet_7_93_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_94_0_clk (.A(clknet_6_47_0_clk),
    .X(clknet_7_94_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_95_0_clk (.A(clknet_6_47_0_clk),
    .X(clknet_7_95_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_96_0_clk (.A(clknet_6_48_0_clk),
    .X(clknet_7_96_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_97_0_clk (.A(clknet_6_48_0_clk),
    .X(clknet_7_97_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_98_0_clk (.A(clknet_6_49_0_clk),
    .X(clknet_7_98_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_99_0_clk (.A(clknet_6_49_0_clk),
    .X(clknet_7_99_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_100_0_clk (.A(clknet_6_50_0_clk),
    .X(clknet_7_100_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_101_0_clk (.A(clknet_6_50_0_clk),
    .X(clknet_7_101_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_102_0_clk (.A(clknet_6_51_0_clk),
    .X(clknet_7_102_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_103_0_clk (.A(clknet_6_51_0_clk),
    .X(clknet_7_103_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_104_0_clk (.A(clknet_6_52_0_clk),
    .X(clknet_7_104_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_105_0_clk (.A(clknet_6_52_0_clk),
    .X(clknet_7_105_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_106_0_clk (.A(clknet_6_53_0_clk),
    .X(clknet_7_106_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_107_0_clk (.A(clknet_6_53_0_clk),
    .X(clknet_7_107_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_108_0_clk (.A(clknet_6_54_0_clk),
    .X(clknet_7_108_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_109_0_clk (.A(clknet_6_54_0_clk),
    .X(clknet_7_109_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_110_0_clk (.A(clknet_6_55_0_clk),
    .X(clknet_7_110_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_111_0_clk (.A(clknet_6_55_0_clk),
    .X(clknet_7_111_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_112_0_clk (.A(clknet_6_56_0_clk),
    .X(clknet_7_112_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_113_0_clk (.A(clknet_6_56_0_clk),
    .X(clknet_7_113_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_114_0_clk (.A(clknet_6_57_0_clk),
    .X(clknet_7_114_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_115_0_clk (.A(clknet_6_57_0_clk),
    .X(clknet_7_115_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_116_0_clk (.A(clknet_6_58_0_clk),
    .X(clknet_7_116_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_117_0_clk (.A(clknet_6_58_0_clk),
    .X(clknet_7_117_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_118_0_clk (.A(clknet_6_59_0_clk),
    .X(clknet_7_118_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_119_0_clk (.A(clknet_6_59_0_clk),
    .X(clknet_7_119_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_120_0_clk (.A(clknet_6_60_0_clk),
    .X(clknet_7_120_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_121_0_clk (.A(clknet_6_60_0_clk),
    .X(clknet_7_121_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_122_0_clk (.A(clknet_6_61_0_clk),
    .X(clknet_7_122_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_123_0_clk (.A(clknet_6_61_0_clk),
    .X(clknet_7_123_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_124_0_clk (.A(clknet_6_62_0_clk),
    .X(clknet_7_124_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_125_0_clk (.A(clknet_6_62_0_clk),
    .X(clknet_7_125_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_126_0_clk (.A(clknet_6_63_0_clk),
    .X(clknet_7_126_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_7_127_0_clk (.A(clknet_6_63_0_clk),
    .X(clknet_7_127_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_0_0_clk (.A(clknet_7_0_0_clk),
    .X(clknet_8_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_1_0_clk (.A(clknet_7_0_0_clk),
    .X(clknet_8_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_2_0_clk (.A(clknet_7_1_0_clk),
    .X(clknet_8_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_3_0_clk (.A(clknet_7_1_0_clk),
    .X(clknet_8_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_4_0_clk (.A(clknet_7_2_0_clk),
    .X(clknet_8_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_5_0_clk (.A(clknet_7_2_0_clk),
    .X(clknet_8_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_6_0_clk (.A(clknet_7_3_0_clk),
    .X(clknet_8_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_7_0_clk (.A(clknet_7_3_0_clk),
    .X(clknet_8_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_8_0_clk (.A(clknet_7_4_0_clk),
    .X(clknet_8_8_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_9_0_clk (.A(clknet_7_4_0_clk),
    .X(clknet_8_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_10_0_clk (.A(clknet_7_5_0_clk),
    .X(clknet_8_10_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_11_0_clk (.A(clknet_7_5_0_clk),
    .X(clknet_8_11_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_12_0_clk (.A(clknet_7_6_0_clk),
    .X(clknet_8_12_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_13_0_clk (.A(clknet_7_6_0_clk),
    .X(clknet_8_13_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_14_0_clk (.A(clknet_7_7_0_clk),
    .X(clknet_8_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_15_0_clk (.A(clknet_7_7_0_clk),
    .X(clknet_8_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_16_0_clk (.A(clknet_7_8_0_clk),
    .X(clknet_8_16_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_17_0_clk (.A(clknet_7_8_0_clk),
    .X(clknet_8_17_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_18_0_clk (.A(clknet_7_9_0_clk),
    .X(clknet_8_18_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_19_0_clk (.A(clknet_7_9_0_clk),
    .X(clknet_8_19_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_20_0_clk (.A(clknet_7_10_0_clk),
    .X(clknet_8_20_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_21_0_clk (.A(clknet_7_10_0_clk),
    .X(clknet_8_21_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_22_0_clk (.A(clknet_7_11_0_clk),
    .X(clknet_8_22_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_23_0_clk (.A(clknet_7_11_0_clk),
    .X(clknet_8_23_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_24_0_clk (.A(clknet_7_12_0_clk),
    .X(clknet_8_24_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_25_0_clk (.A(clknet_7_12_0_clk),
    .X(clknet_8_25_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_26_0_clk (.A(clknet_7_13_0_clk),
    .X(clknet_8_26_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_27_0_clk (.A(clknet_7_13_0_clk),
    .X(clknet_8_27_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_28_0_clk (.A(clknet_7_14_0_clk),
    .X(clknet_8_28_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_29_0_clk (.A(clknet_7_14_0_clk),
    .X(clknet_8_29_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_30_0_clk (.A(clknet_7_15_0_clk),
    .X(clknet_8_30_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_31_0_clk (.A(clknet_7_15_0_clk),
    .X(clknet_8_31_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_32_0_clk (.A(clknet_7_16_0_clk),
    .X(clknet_8_32_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_33_0_clk (.A(clknet_7_16_0_clk),
    .X(clknet_8_33_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_34_0_clk (.A(clknet_7_17_0_clk),
    .X(clknet_8_34_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_35_0_clk (.A(clknet_7_17_0_clk),
    .X(clknet_8_35_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_36_0_clk (.A(clknet_7_18_0_clk),
    .X(clknet_8_36_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_37_0_clk (.A(clknet_7_18_0_clk),
    .X(clknet_8_37_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_38_0_clk (.A(clknet_7_19_0_clk),
    .X(clknet_8_38_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_39_0_clk (.A(clknet_7_19_0_clk),
    .X(clknet_8_39_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_40_0_clk (.A(clknet_7_20_0_clk),
    .X(clknet_8_40_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_41_0_clk (.A(clknet_7_20_0_clk),
    .X(clknet_8_41_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_42_0_clk (.A(clknet_7_21_0_clk),
    .X(clknet_8_42_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_43_0_clk (.A(clknet_7_21_0_clk),
    .X(clknet_8_43_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_44_0_clk (.A(clknet_7_22_0_clk),
    .X(clknet_8_44_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_45_0_clk (.A(clknet_7_22_0_clk),
    .X(clknet_8_45_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_46_0_clk (.A(clknet_7_23_0_clk),
    .X(clknet_8_46_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_47_0_clk (.A(clknet_7_23_0_clk),
    .X(clknet_8_47_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_48_0_clk (.A(clknet_7_24_0_clk),
    .X(clknet_8_48_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_49_0_clk (.A(clknet_7_24_0_clk),
    .X(clknet_8_49_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_50_0_clk (.A(clknet_7_25_0_clk),
    .X(clknet_8_50_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_51_0_clk (.A(clknet_7_25_0_clk),
    .X(clknet_8_51_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_52_0_clk (.A(clknet_7_26_0_clk),
    .X(clknet_8_52_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_53_0_clk (.A(clknet_7_26_0_clk),
    .X(clknet_8_53_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_54_0_clk (.A(clknet_7_27_0_clk),
    .X(clknet_8_54_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_55_0_clk (.A(clknet_7_27_0_clk),
    .X(clknet_8_55_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_56_0_clk (.A(clknet_7_28_0_clk),
    .X(clknet_8_56_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_57_0_clk (.A(clknet_7_28_0_clk),
    .X(clknet_8_57_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_58_0_clk (.A(clknet_7_29_0_clk),
    .X(clknet_8_58_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_59_0_clk (.A(clknet_7_29_0_clk),
    .X(clknet_8_59_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_60_0_clk (.A(clknet_7_30_0_clk),
    .X(clknet_8_60_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_61_0_clk (.A(clknet_7_30_0_clk),
    .X(clknet_8_61_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_62_0_clk (.A(clknet_7_31_0_clk),
    .X(clknet_8_62_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_63_0_clk (.A(clknet_7_31_0_clk),
    .X(clknet_8_63_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_64_0_clk (.A(clknet_7_32_0_clk),
    .X(clknet_8_64_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_65_0_clk (.A(clknet_7_32_0_clk),
    .X(clknet_8_65_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_66_0_clk (.A(clknet_7_33_0_clk),
    .X(clknet_8_66_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_67_0_clk (.A(clknet_7_33_0_clk),
    .X(clknet_8_67_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_68_0_clk (.A(clknet_7_34_0_clk),
    .X(clknet_8_68_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_69_0_clk (.A(clknet_7_34_0_clk),
    .X(clknet_8_69_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_70_0_clk (.A(clknet_7_35_0_clk),
    .X(clknet_8_70_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_71_0_clk (.A(clknet_7_35_0_clk),
    .X(clknet_8_71_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_72_0_clk (.A(clknet_7_36_0_clk),
    .X(clknet_8_72_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_73_0_clk (.A(clknet_7_36_0_clk),
    .X(clknet_8_73_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_74_0_clk (.A(clknet_7_37_0_clk),
    .X(clknet_8_74_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_75_0_clk (.A(clknet_7_37_0_clk),
    .X(clknet_8_75_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_76_0_clk (.A(clknet_7_38_0_clk),
    .X(clknet_8_76_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_77_0_clk (.A(clknet_7_38_0_clk),
    .X(clknet_8_77_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_78_0_clk (.A(clknet_7_39_0_clk),
    .X(clknet_8_78_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_79_0_clk (.A(clknet_7_39_0_clk),
    .X(clknet_8_79_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_80_0_clk (.A(clknet_7_40_0_clk),
    .X(clknet_8_80_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_81_0_clk (.A(clknet_7_40_0_clk),
    .X(clknet_8_81_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_82_0_clk (.A(clknet_7_41_0_clk),
    .X(clknet_8_82_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_83_0_clk (.A(clknet_7_41_0_clk),
    .X(clknet_8_83_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_84_0_clk (.A(clknet_7_42_0_clk),
    .X(clknet_8_84_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_85_0_clk (.A(clknet_7_42_0_clk),
    .X(clknet_8_85_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_86_0_clk (.A(clknet_7_43_0_clk),
    .X(clknet_8_86_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_87_0_clk (.A(clknet_7_43_0_clk),
    .X(clknet_8_87_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_88_0_clk (.A(clknet_7_44_0_clk),
    .X(clknet_8_88_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_89_0_clk (.A(clknet_7_44_0_clk),
    .X(clknet_8_89_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_90_0_clk (.A(clknet_7_45_0_clk),
    .X(clknet_8_90_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_91_0_clk (.A(clknet_7_45_0_clk),
    .X(clknet_8_91_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_92_0_clk (.A(clknet_7_46_0_clk),
    .X(clknet_8_92_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_93_0_clk (.A(clknet_7_46_0_clk),
    .X(clknet_8_93_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_94_0_clk (.A(clknet_7_47_0_clk),
    .X(clknet_8_94_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_95_0_clk (.A(clknet_7_47_0_clk),
    .X(clknet_8_95_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_96_0_clk (.A(clknet_7_48_0_clk),
    .X(clknet_8_96_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_97_0_clk (.A(clknet_7_48_0_clk),
    .X(clknet_8_97_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_98_0_clk (.A(clknet_7_49_0_clk),
    .X(clknet_8_98_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_99_0_clk (.A(clknet_7_49_0_clk),
    .X(clknet_8_99_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_100_0_clk (.A(clknet_7_50_0_clk),
    .X(clknet_8_100_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_101_0_clk (.A(clknet_7_50_0_clk),
    .X(clknet_8_101_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_102_0_clk (.A(clknet_7_51_0_clk),
    .X(clknet_8_102_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_103_0_clk (.A(clknet_7_51_0_clk),
    .X(clknet_8_103_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_104_0_clk (.A(clknet_7_52_0_clk),
    .X(clknet_8_104_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_105_0_clk (.A(clknet_7_52_0_clk),
    .X(clknet_8_105_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_106_0_clk (.A(clknet_7_53_0_clk),
    .X(clknet_8_106_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_107_0_clk (.A(clknet_7_53_0_clk),
    .X(clknet_8_107_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_108_0_clk (.A(clknet_7_54_0_clk),
    .X(clknet_8_108_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_109_0_clk (.A(clknet_7_54_0_clk),
    .X(clknet_8_109_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_110_0_clk (.A(clknet_7_55_0_clk),
    .X(clknet_8_110_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_111_0_clk (.A(clknet_7_55_0_clk),
    .X(clknet_8_111_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_112_0_clk (.A(clknet_7_56_0_clk),
    .X(clknet_8_112_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_113_0_clk (.A(clknet_7_56_0_clk),
    .X(clknet_8_113_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_114_0_clk (.A(clknet_7_57_0_clk),
    .X(clknet_8_114_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_115_0_clk (.A(clknet_7_57_0_clk),
    .X(clknet_8_115_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_116_0_clk (.A(clknet_7_58_0_clk),
    .X(clknet_8_116_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_117_0_clk (.A(clknet_7_58_0_clk),
    .X(clknet_8_117_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_118_0_clk (.A(clknet_7_59_0_clk),
    .X(clknet_8_118_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_119_0_clk (.A(clknet_7_59_0_clk),
    .X(clknet_8_119_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_120_0_clk (.A(clknet_7_60_0_clk),
    .X(clknet_8_120_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_121_0_clk (.A(clknet_7_60_0_clk),
    .X(clknet_8_121_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_122_0_clk (.A(clknet_7_61_0_clk),
    .X(clknet_8_122_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_123_0_clk (.A(clknet_7_61_0_clk),
    .X(clknet_8_123_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_124_0_clk (.A(clknet_7_62_0_clk),
    .X(clknet_8_124_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_125_0_clk (.A(clknet_7_62_0_clk),
    .X(clknet_8_125_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_126_0_clk (.A(clknet_7_63_0_clk),
    .X(clknet_8_126_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_127_0_clk (.A(clknet_7_63_0_clk),
    .X(clknet_8_127_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_128_0_clk (.A(clknet_7_64_0_clk),
    .X(clknet_8_128_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_129_0_clk (.A(clknet_7_64_0_clk),
    .X(clknet_8_129_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_130_0_clk (.A(clknet_7_65_0_clk),
    .X(clknet_8_130_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_131_0_clk (.A(clknet_7_65_0_clk),
    .X(clknet_8_131_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_132_0_clk (.A(clknet_7_66_0_clk),
    .X(clknet_8_132_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_133_0_clk (.A(clknet_7_66_0_clk),
    .X(clknet_8_133_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_134_0_clk (.A(clknet_7_67_0_clk),
    .X(clknet_8_134_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_135_0_clk (.A(clknet_7_67_0_clk),
    .X(clknet_8_135_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_136_0_clk (.A(clknet_7_68_0_clk),
    .X(clknet_8_136_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_137_0_clk (.A(clknet_7_68_0_clk),
    .X(clknet_8_137_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_138_0_clk (.A(clknet_7_69_0_clk),
    .X(clknet_8_138_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_139_0_clk (.A(clknet_7_69_0_clk),
    .X(clknet_8_139_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_140_0_clk (.A(clknet_7_70_0_clk),
    .X(clknet_8_140_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_141_0_clk (.A(clknet_7_70_0_clk),
    .X(clknet_8_141_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_142_0_clk (.A(clknet_7_71_0_clk),
    .X(clknet_8_142_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_143_0_clk (.A(clknet_7_71_0_clk),
    .X(clknet_8_143_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_144_0_clk (.A(clknet_7_72_0_clk),
    .X(clknet_8_144_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_145_0_clk (.A(clknet_7_72_0_clk),
    .X(clknet_8_145_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_146_0_clk (.A(clknet_7_73_0_clk),
    .X(clknet_8_146_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_147_0_clk (.A(clknet_7_73_0_clk),
    .X(clknet_8_147_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_148_0_clk (.A(clknet_7_74_0_clk),
    .X(clknet_8_148_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_149_0_clk (.A(clknet_7_74_0_clk),
    .X(clknet_8_149_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_150_0_clk (.A(clknet_7_75_0_clk),
    .X(clknet_8_150_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_151_0_clk (.A(clknet_7_75_0_clk),
    .X(clknet_8_151_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_152_0_clk (.A(clknet_7_76_0_clk),
    .X(clknet_8_152_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_153_0_clk (.A(clknet_7_76_0_clk),
    .X(clknet_8_153_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_154_0_clk (.A(clknet_7_77_0_clk),
    .X(clknet_8_154_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_155_0_clk (.A(clknet_7_77_0_clk),
    .X(clknet_8_155_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_156_0_clk (.A(clknet_7_78_0_clk),
    .X(clknet_8_156_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_157_0_clk (.A(clknet_7_78_0_clk),
    .X(clknet_8_157_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_158_0_clk (.A(clknet_7_79_0_clk),
    .X(clknet_8_158_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_159_0_clk (.A(clknet_7_79_0_clk),
    .X(clknet_8_159_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_160_0_clk (.A(clknet_7_80_0_clk),
    .X(clknet_8_160_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_161_0_clk (.A(clknet_7_80_0_clk),
    .X(clknet_8_161_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_162_0_clk (.A(clknet_7_81_0_clk),
    .X(clknet_8_162_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_163_0_clk (.A(clknet_7_81_0_clk),
    .X(clknet_8_163_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_164_0_clk (.A(clknet_7_82_0_clk),
    .X(clknet_8_164_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_165_0_clk (.A(clknet_7_82_0_clk),
    .X(clknet_8_165_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_166_0_clk (.A(clknet_7_83_0_clk),
    .X(clknet_8_166_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_167_0_clk (.A(clknet_7_83_0_clk),
    .X(clknet_8_167_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_168_0_clk (.A(clknet_7_84_0_clk),
    .X(clknet_8_168_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_169_0_clk (.A(clknet_7_84_0_clk),
    .X(clknet_8_169_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_170_0_clk (.A(clknet_7_85_0_clk),
    .X(clknet_8_170_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_171_0_clk (.A(clknet_7_85_0_clk),
    .X(clknet_8_171_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_172_0_clk (.A(clknet_7_86_0_clk),
    .X(clknet_8_172_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_173_0_clk (.A(clknet_7_86_0_clk),
    .X(clknet_8_173_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_174_0_clk (.A(clknet_7_87_0_clk),
    .X(clknet_8_174_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_175_0_clk (.A(clknet_7_87_0_clk),
    .X(clknet_8_175_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_176_0_clk (.A(clknet_7_88_0_clk),
    .X(clknet_8_176_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_177_0_clk (.A(clknet_7_88_0_clk),
    .X(clknet_8_177_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_178_0_clk (.A(clknet_7_89_0_clk),
    .X(clknet_8_178_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_179_0_clk (.A(clknet_7_89_0_clk),
    .X(clknet_8_179_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_180_0_clk (.A(clknet_7_90_0_clk),
    .X(clknet_8_180_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_181_0_clk (.A(clknet_7_90_0_clk),
    .X(clknet_8_181_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_182_0_clk (.A(clknet_7_91_0_clk),
    .X(clknet_8_182_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_183_0_clk (.A(clknet_7_91_0_clk),
    .X(clknet_8_183_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_184_0_clk (.A(clknet_7_92_0_clk),
    .X(clknet_8_184_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_185_0_clk (.A(clknet_7_92_0_clk),
    .X(clknet_8_185_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_186_0_clk (.A(clknet_7_93_0_clk),
    .X(clknet_8_186_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_187_0_clk (.A(clknet_7_93_0_clk),
    .X(clknet_8_187_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_188_0_clk (.A(clknet_7_94_0_clk),
    .X(clknet_8_188_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_189_0_clk (.A(clknet_7_94_0_clk),
    .X(clknet_8_189_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_190_0_clk (.A(clknet_7_95_0_clk),
    .X(clknet_8_190_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_191_0_clk (.A(clknet_7_95_0_clk),
    .X(clknet_8_191_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_192_0_clk (.A(clknet_7_96_0_clk),
    .X(clknet_8_192_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_193_0_clk (.A(clknet_7_96_0_clk),
    .X(clknet_8_193_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_194_0_clk (.A(clknet_7_97_0_clk),
    .X(clknet_8_194_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_195_0_clk (.A(clknet_7_97_0_clk),
    .X(clknet_8_195_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_196_0_clk (.A(clknet_7_98_0_clk),
    .X(clknet_8_196_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_197_0_clk (.A(clknet_7_98_0_clk),
    .X(clknet_8_197_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_198_0_clk (.A(clknet_7_99_0_clk),
    .X(clknet_8_198_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_199_0_clk (.A(clknet_7_99_0_clk),
    .X(clknet_8_199_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_200_0_clk (.A(clknet_7_100_0_clk),
    .X(clknet_8_200_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_201_0_clk (.A(clknet_7_100_0_clk),
    .X(clknet_8_201_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_202_0_clk (.A(clknet_7_101_0_clk),
    .X(clknet_8_202_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_203_0_clk (.A(clknet_7_101_0_clk),
    .X(clknet_8_203_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_204_0_clk (.A(clknet_7_102_0_clk),
    .X(clknet_8_204_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_205_0_clk (.A(clknet_7_102_0_clk),
    .X(clknet_8_205_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_206_0_clk (.A(clknet_7_103_0_clk),
    .X(clknet_8_206_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_207_0_clk (.A(clknet_7_103_0_clk),
    .X(clknet_8_207_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_208_0_clk (.A(clknet_7_104_0_clk),
    .X(clknet_8_208_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_209_0_clk (.A(clknet_7_104_0_clk),
    .X(clknet_8_209_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_210_0_clk (.A(clknet_7_105_0_clk),
    .X(clknet_8_210_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_211_0_clk (.A(clknet_7_105_0_clk),
    .X(clknet_8_211_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_212_0_clk (.A(clknet_7_106_0_clk),
    .X(clknet_8_212_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_213_0_clk (.A(clknet_7_106_0_clk),
    .X(clknet_8_213_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_214_0_clk (.A(clknet_7_107_0_clk),
    .X(clknet_8_214_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_215_0_clk (.A(clknet_7_107_0_clk),
    .X(clknet_8_215_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_216_0_clk (.A(clknet_7_108_0_clk),
    .X(clknet_8_216_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_217_0_clk (.A(clknet_7_108_0_clk),
    .X(clknet_8_217_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_218_0_clk (.A(clknet_7_109_0_clk),
    .X(clknet_8_218_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_219_0_clk (.A(clknet_7_109_0_clk),
    .X(clknet_8_219_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_220_0_clk (.A(clknet_7_110_0_clk),
    .X(clknet_8_220_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_221_0_clk (.A(clknet_7_110_0_clk),
    .X(clknet_8_221_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_222_0_clk (.A(clknet_7_111_0_clk),
    .X(clknet_8_222_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_223_0_clk (.A(clknet_7_111_0_clk),
    .X(clknet_8_223_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_224_0_clk (.A(clknet_7_112_0_clk),
    .X(clknet_8_224_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_225_0_clk (.A(clknet_7_112_0_clk),
    .X(clknet_8_225_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_226_0_clk (.A(clknet_7_113_0_clk),
    .X(clknet_8_226_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_227_0_clk (.A(clknet_7_113_0_clk),
    .X(clknet_8_227_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_228_0_clk (.A(clknet_7_114_0_clk),
    .X(clknet_8_228_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_229_0_clk (.A(clknet_7_114_0_clk),
    .X(clknet_8_229_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_230_0_clk (.A(clknet_7_115_0_clk),
    .X(clknet_8_230_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_231_0_clk (.A(clknet_7_115_0_clk),
    .X(clknet_8_231_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_232_0_clk (.A(clknet_7_116_0_clk),
    .X(clknet_8_232_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_233_0_clk (.A(clknet_7_116_0_clk),
    .X(clknet_8_233_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_234_0_clk (.A(clknet_7_117_0_clk),
    .X(clknet_8_234_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_235_0_clk (.A(clknet_7_117_0_clk),
    .X(clknet_8_235_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_236_0_clk (.A(clknet_7_118_0_clk),
    .X(clknet_8_236_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_237_0_clk (.A(clknet_7_118_0_clk),
    .X(clknet_8_237_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_238_0_clk (.A(clknet_7_119_0_clk),
    .X(clknet_8_238_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_239_0_clk (.A(clknet_7_119_0_clk),
    .X(clknet_8_239_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_240_0_clk (.A(clknet_7_120_0_clk),
    .X(clknet_8_240_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_241_0_clk (.A(clknet_7_120_0_clk),
    .X(clknet_8_241_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_242_0_clk (.A(clknet_7_121_0_clk),
    .X(clknet_8_242_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_243_0_clk (.A(clknet_7_121_0_clk),
    .X(clknet_8_243_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_244_0_clk (.A(clknet_7_122_0_clk),
    .X(clknet_8_244_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_245_0_clk (.A(clknet_7_122_0_clk),
    .X(clknet_8_245_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_246_0_clk (.A(clknet_7_123_0_clk),
    .X(clknet_8_246_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_247_0_clk (.A(clknet_7_123_0_clk),
    .X(clknet_8_247_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_248_0_clk (.A(clknet_7_124_0_clk),
    .X(clknet_8_248_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_249_0_clk (.A(clknet_7_124_0_clk),
    .X(clknet_8_249_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_250_0_clk (.A(clknet_7_125_0_clk),
    .X(clknet_8_250_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_251_0_clk (.A(clknet_7_125_0_clk),
    .X(clknet_8_251_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_252_0_clk (.A(clknet_7_126_0_clk),
    .X(clknet_8_252_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_253_0_clk (.A(clknet_7_126_0_clk),
    .X(clknet_8_253_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_254_0_clk (.A(clknet_7_127_0_clk),
    .X(clknet_8_254_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_8_255_0_clk (.A(clknet_7_127_0_clk),
    .X(clknet_8_255_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_clk (.A(clknet_8_255_0_clk),
    .X(clknet_opt_0_clk));
endmodule
