`ifndef SP_DEFAULT
`define SP_DEFAULT
/*
Copyright (c) 2015, Steven F. Hoover

Redistribution and use in source and binary forms, with or without
modification, are permitted provided that the following conditions are met:

    * Redistributions of source code must retain the above copyright notice,
      this list of conditions and the following disclaimer.
    * Redistributions in binary form must reproduce the above copyright
      notice, this list of conditions and the following disclaimer in the
      documentation and/or other materials provided with the distribution.
    * The name of Steven F. Hoover
      may not be used to endorse or promote products derived from this software
      without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE
FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/


// File included by SandPiper-generated code for the default project configuration.
`include "includes/sandpiper.vh"


// Latch macros.  Inject 'x in simulation for clk === 'x.

// A-phase latch.
`ifdef SP_PHYS
`define TLV_LATCH(in, out, clk) \
always @ (in, clk) begin        \
  if (clk === 1'b1)             \
    out <= in;                  \
  else if (clk === 1'bx)        \
    out <= 'x;                  \
end
`else
`define TLV_LATCH(in, out, clk) always @ (in, clk) if (clk == 1'b1) out <= in;
`endif  // SP_PHYS

// B-phase latch.
`ifdef SP_PHYS
`define TLV_BLATCH(out, in, clk) \
always @ (in, clk) begin         \
  if (!clk === 1'b1)             \
    out <= in;                   \
  else if (!clk === 1'bx)        \
    out <= 'x;                   \
end
`else
`define TLV_BLATCH(out, in, clk) always @ (in, clk) if (!clk == 1'b1) out <= in;
`endif  // SP_PHYS


	   
`endif  // SP_DEFAULT
